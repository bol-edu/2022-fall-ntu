
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "pp_loop_interface.svh"
`include "pp_loop_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_dpu_keygen.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_dpu_keygen.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_dpu_keygen.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_read_p2_fu_664.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_read_p2_fu_664.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_read_p2_fu_664.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.grp_read_p1_fu_165.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.grp_read_p1_fu_165.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.grp_read_p1_fu_165.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.call_ln290_write_p3_fu_181.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.call_ln290_write_p3_fu_181.ap_ready;
    assign module_intf_6.ap_done = 1'b0;
    assign module_intf_6.ap_continue = 1'b0;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.call_ln291_write_p4_fu_189.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.call_ln291_write_p4_fu_189.ap_ready;
    assign module_intf_7.ap_done = 1'b0;
    assign module_intf_7.ap_continue = 1'b0;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.grp_read_p1_fu_145.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.grp_read_p1_fu_145.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.grp_read_p1_fu_145.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.call_ln281_write_p3_fu_161.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.call_ln281_write_p3_fu_161.ap_ready;
    assign module_intf_10.ap_done = 1'b0;
    assign module_intf_10.ap_continue = 1'b0;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.grp_read_p1_fu_155.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.grp_read_p1_fu_155.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.grp_read_p1_fu_155.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.grp_read_p2_fu_162.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.grp_read_p2_fu_162.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.grp_read_p2_fu_162.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.call_ln193_write_p3_fu_178.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.call_ln193_write_p3_fu_178.ap_ready;
    assign module_intf_14.ap_done = 1'b0;
    assign module_intf_14.ap_continue = 1'b0;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.call_ln194_write_p4_fu_186.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.call_ln194_write_p4_fu_186.ap_ready;
    assign module_intf_15.ap_done = 1'b0;
    assign module_intf_15.ap_continue = 1'b0;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.grp_read_p1_fu_147.ap_start;
    assign module_intf_17.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.grp_read_p1_fu_147.ap_ready;
    assign module_intf_17.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.grp_read_p1_fu_147.ap_done;
    assign module_intf_17.ap_continue = 1'b1;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.call_ln164_write_p3_fu_163.ap_start;
    assign module_intf_18.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.call_ln164_write_p3_fu_163.ap_ready;
    assign module_intf_18.ap_done = 1'b0;
    assign module_intf_18.ap_continue = 1'b0;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.grp_read_p1_fu_178.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.grp_read_p1_fu_178.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.grp_read_p1_fu_178.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.grp_read_p2_fu_185.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.grp_read_p2_fu_185.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.grp_read_p2_fu_185.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = 1'b0;
    assign module_intf_22.ap_ready = 1'b0;
    assign module_intf_22.ap_done = 1'b0;
    assign module_intf_22.ap_continue = 1'b0;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.call_ln154_write_p3_fu_201.ap_start;
    assign module_intf_23.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.call_ln154_write_p3_fu_201.ap_ready;
    assign module_intf_23.ap_done = 1'b0;
    assign module_intf_23.ap_continue = 1'b0;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.grp_read_p1_fu_178.ap_start;
    assign module_intf_25.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.grp_read_p1_fu_178.ap_ready;
    assign module_intf_25.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.grp_read_p1_fu_178.ap_done;
    assign module_intf_25.ap_continue = 1'b1;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.grp_read_p2_fu_185.ap_start;
    assign module_intf_26.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.grp_read_p2_fu_185.ap_ready;
    assign module_intf_26.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.grp_read_p2_fu_185.ap_done;
    assign module_intf_26.ap_continue = 1'b1;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.call_ln144_write_p3_fu_201.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.call_ln144_write_p3_fu_201.ap_ready;
    assign module_intf_27.ap_done = 1'b0;
    assign module_intf_27.ap_continue = 1'b0;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_start;
    assign module_intf_28.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_ready;
    assign module_intf_28.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_done;
    assign module_intf_28.ap_continue = 1'b1;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.grp_read_p1_fu_151.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.grp_read_p1_fu_151.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.grp_read_p1_fu_151.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.call_ln302_write_p3_fu_167.ap_start;
    assign module_intf_30.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.call_ln302_write_p3_fu_167.ap_ready;
    assign module_intf_30.ap_done = 1'b0;
    assign module_intf_30.ap_continue = 1'b0;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.call_ln303_write_p4_fu_175.ap_start;
    assign module_intf_31.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.call_ln303_write_p4_fu_175.ap_ready;
    assign module_intf_31.ap_done = 1'b0;
    assign module_intf_31.ap_continue = 1'b0;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.grp_read_p1_fu_137.ap_start;
    assign module_intf_33.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.grp_read_p1_fu_137.ap_ready;
    assign module_intf_33.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.grp_read_p1_fu_137.ap_done;
    assign module_intf_33.ap_continue = 1'b1;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.call_ln312_write_p3_fu_153.ap_start;
    assign module_intf_34.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.call_ln312_write_p3_fu_153.ap_ready;
    assign module_intf_34.ap_done = 1'b0;
    assign module_intf_34.ap_continue = 1'b0;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_start;
    assign module_intf_35.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_ready;
    assign module_intf_35.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_done;
    assign module_intf_35.ap_continue = 1'b1;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.grp_read_p1_fu_137.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.grp_read_p1_fu_137.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.grp_read_p1_fu_137.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.call_ln321_write_p4_fu_153.ap_start;
    assign module_intf_37.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.call_ln321_write_p4_fu_153.ap_ready;
    assign module_intf_37.ap_done = 1'b0;
    assign module_intf_37.ap_continue = 1'b0;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_start;
    assign module_intf_38.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_ready;
    assign module_intf_38.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_done;
    assign module_intf_38.ap_continue = 1'b1;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.grp_read_p1_fu_164.ap_start;
    assign module_intf_39.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.grp_read_p1_fu_164.ap_ready;
    assign module_intf_39.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.grp_read_p1_fu_164.ap_done;
    assign module_intf_39.ap_continue = 1'b1;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.grp_read_p2_fu_171.ap_start;
    assign module_intf_40.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.grp_read_p2_fu_171.ap_ready;
    assign module_intf_40.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.grp_read_p2_fu_171.ap_done;
    assign module_intf_40.ap_continue = 1'b1;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.call_ln330_write_p3_fu_187.ap_start;
    assign module_intf_41.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.call_ln330_write_p3_fu_187.ap_ready;
    assign module_intf_41.ap_done = 1'b0;
    assign module_intf_41.ap_continue = 1'b0;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_start;
    assign module_intf_42.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_ready;
    assign module_intf_42.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_done;
    assign module_intf_42.ap_continue = 1'b1;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.grp_read_ntt_fu_112.ap_start;
    assign module_intf_43.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.grp_read_ntt_fu_112.ap_ready;
    assign module_intf_43.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.grp_read_ntt_fu_112.ap_done;
    assign module_intf_43.ap_continue = 1'b1;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.call_ln338_write_p3_fu_128.ap_start;
    assign module_intf_44.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.call_ln338_write_p3_fu_128.ap_ready;
    assign module_intf_44.ap_done = 1'b0;
    assign module_intf_44.ap_continue = 1'b0;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_start;
    assign module_intf_45.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_ready;
    assign module_intf_45.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_done;
    assign module_intf_45.ap_continue = 1'b1;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.grp_read_p1_fu_165.ap_start;
    assign module_intf_46.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.grp_read_p1_fu_165.ap_ready;
    assign module_intf_46.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.grp_read_p1_fu_165.ap_done;
    assign module_intf_46.ap_continue = 1'b1;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.grp_read_p2_fu_172.ap_start;
    assign module_intf_47.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.grp_read_p2_fu_172.ap_ready;
    assign module_intf_47.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.grp_read_p2_fu_172.ap_done;
    assign module_intf_47.ap_continue = 1'b1;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.call_ln233_write_p3_fu_188.ap_start;
    assign module_intf_48.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.call_ln233_write_p3_fu_188.ap_ready;
    assign module_intf_48.ap_done = 1'b0;
    assign module_intf_48.ap_continue = 1'b0;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.call_ln234_write_p4_fu_196.ap_start;
    assign module_intf_49.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.call_ln234_write_p4_fu_196.ap_ready;
    assign module_intf_49.ap_done = 1'b0;
    assign module_intf_49.ap_continue = 1'b0;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_start;
    assign module_intf_50.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_ready;
    assign module_intf_50.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_done;
    assign module_intf_50.ap_continue = 1'b1;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.grp_read_p1_fu_137.ap_start;
    assign module_intf_51.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.grp_read_p1_fu_137.ap_ready;
    assign module_intf_51.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.grp_read_p1_fu_137.ap_done;
    assign module_intf_51.ap_continue = 1'b1;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.call_ln243_write_p3_fu_153.ap_start;
    assign module_intf_52.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.call_ln243_write_p3_fu_153.ap_ready;
    assign module_intf_52.ap_done = 1'b0;
    assign module_intf_52.ap_continue = 1'b0;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;
    nodf_module_intf module_intf_53(clock,reset);
    assign module_intf_53.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_start;
    assign module_intf_53.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_ready;
    assign module_intf_53.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_done;
    assign module_intf_53.ap_continue = 1'b1;
    assign module_intf_53.finish = finish;
    csv_file_dump mstatus_csv_dumper_53;
    nodf_module_monitor module_monitor_53;
    nodf_module_intf module_intf_54(clock,reset);
    assign module_intf_54.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.grp_read_p1_fu_137.ap_start;
    assign module_intf_54.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.grp_read_p1_fu_137.ap_ready;
    assign module_intf_54.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.grp_read_p1_fu_137.ap_done;
    assign module_intf_54.ap_continue = 1'b1;
    assign module_intf_54.finish = finish;
    csv_file_dump mstatus_csv_dumper_54;
    nodf_module_monitor module_monitor_54;
    nodf_module_intf module_intf_55(clock,reset);
    assign module_intf_55.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.call_ln252_write_p4_fu_153.ap_start;
    assign module_intf_55.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.call_ln252_write_p4_fu_153.ap_ready;
    assign module_intf_55.ap_done = 1'b0;
    assign module_intf_55.ap_continue = 1'b0;
    assign module_intf_55.finish = finish;
    csv_file_dump mstatus_csv_dumper_55;
    nodf_module_monitor module_monitor_55;
    nodf_module_intf module_intf_56(clock,reset);
    assign module_intf_56.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_start;
    assign module_intf_56.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_ready;
    assign module_intf_56.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_done;
    assign module_intf_56.ap_continue = 1'b1;
    assign module_intf_56.finish = finish;
    csv_file_dump mstatus_csv_dumper_56;
    nodf_module_monitor module_monitor_56;
    nodf_module_intf module_intf_57(clock,reset);
    assign module_intf_57.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.grp_read_p1_fu_154.ap_start;
    assign module_intf_57.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.grp_read_p1_fu_154.ap_ready;
    assign module_intf_57.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.grp_read_p1_fu_154.ap_done;
    assign module_intf_57.ap_continue = 1'b1;
    assign module_intf_57.finish = finish;
    csv_file_dump mstatus_csv_dumper_57;
    nodf_module_monitor module_monitor_57;
    nodf_module_intf module_intf_58(clock,reset);
    assign module_intf_58.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.grp_read_p2_fu_161.ap_start;
    assign module_intf_58.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.grp_read_p2_fu_161.ap_ready;
    assign module_intf_58.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.grp_read_p2_fu_161.ap_done;
    assign module_intf_58.ap_continue = 1'b1;
    assign module_intf_58.finish = finish;
    csv_file_dump mstatus_csv_dumper_58;
    nodf_module_monitor module_monitor_58;
    nodf_module_intf module_intf_59(clock,reset);
    assign module_intf_59.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.call_ln261_write_p3_fu_177.ap_start;
    assign module_intf_59.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.call_ln261_write_p3_fu_177.ap_ready;
    assign module_intf_59.ap_done = 1'b0;
    assign module_intf_59.ap_continue = 1'b0;
    assign module_intf_59.finish = finish;
    csv_file_dump mstatus_csv_dumper_59;
    nodf_module_monitor module_monitor_59;
    nodf_module_intf module_intf_60(clock,reset);
    assign module_intf_60.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_start;
    assign module_intf_60.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_ready;
    assign module_intf_60.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_done;
    assign module_intf_60.ap_continue = 1'b1;
    assign module_intf_60.finish = finish;
    csv_file_dump mstatus_csv_dumper_60;
    nodf_module_monitor module_monitor_60;
    nodf_module_intf module_intf_61(clock,reset);
    assign module_intf_61.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.grp_read_p1_fu_127.ap_start;
    assign module_intf_61.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.grp_read_p1_fu_127.ap_ready;
    assign module_intf_61.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.grp_read_p1_fu_127.ap_done;
    assign module_intf_61.ap_continue = 1'b1;
    assign module_intf_61.finish = finish;
    csv_file_dump mstatus_csv_dumper_61;
    nodf_module_monitor module_monitor_61;
    nodf_module_intf module_intf_62(clock,reset);
    assign module_intf_62.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.grp_read_p2_fu_134.ap_start;
    assign module_intf_62.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.grp_read_p2_fu_134.ap_ready;
    assign module_intf_62.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.grp_read_p2_fu_134.ap_done;
    assign module_intf_62.ap_continue = 1'b1;
    assign module_intf_62.finish = finish;
    csv_file_dump mstatus_csv_dumper_62;
    nodf_module_monitor module_monitor_62;
    nodf_module_intf module_intf_63(clock,reset);
    assign module_intf_63.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.call_ln271_write_p3_fu_151.ap_start;
    assign module_intf_63.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.call_ln271_write_p3_fu_151.ap_ready;
    assign module_intf_63.ap_done = 1'b0;
    assign module_intf_63.ap_continue = 1'b0;
    assign module_intf_63.finish = finish;
    csv_file_dump mstatus_csv_dumper_63;
    nodf_module_monitor module_monitor_63;
    nodf_module_intf module_intf_64(clock,reset);
    assign module_intf_64.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_start;
    assign module_intf_64.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_ready;
    assign module_intf_64.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_done;
    assign module_intf_64.ap_continue = 1'b1;
    assign module_intf_64.finish = finish;
    csv_file_dump mstatus_csv_dumper_64;
    nodf_module_monitor module_monitor_64;
    nodf_module_intf module_intf_65(clock,reset);
    assign module_intf_65.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.grp_read_p1_fu_137.ap_start;
    assign module_intf_65.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.grp_read_p1_fu_137.ap_ready;
    assign module_intf_65.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.grp_read_p1_fu_137.ap_done;
    assign module_intf_65.ap_continue = 1'b1;
    assign module_intf_65.finish = finish;
    csv_file_dump mstatus_csv_dumper_65;
    nodf_module_monitor module_monitor_65;
    nodf_module_intf module_intf_66(clock,reset);
    assign module_intf_66.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.call_ln203_write_p3_fu_153.ap_start;
    assign module_intf_66.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.call_ln203_write_p3_fu_153.ap_ready;
    assign module_intf_66.ap_done = 1'b0;
    assign module_intf_66.ap_continue = 1'b0;
    assign module_intf_66.finish = finish;
    csv_file_dump mstatus_csv_dumper_66;
    nodf_module_monitor module_monitor_66;
    nodf_module_intf module_intf_67(clock,reset);
    assign module_intf_67.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_start;
    assign module_intf_67.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_ready;
    assign module_intf_67.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_done;
    assign module_intf_67.ap_continue = 1'b1;
    assign module_intf_67.finish = finish;
    csv_file_dump mstatus_csv_dumper_67;
    nodf_module_monitor module_monitor_67;
    nodf_module_intf module_intf_68(clock,reset);
    assign module_intf_68.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.grp_read_p1_fu_137.ap_start;
    assign module_intf_68.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.grp_read_p1_fu_137.ap_ready;
    assign module_intf_68.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.grp_read_p1_fu_137.ap_done;
    assign module_intf_68.ap_continue = 1'b1;
    assign module_intf_68.finish = finish;
    csv_file_dump mstatus_csv_dumper_68;
    nodf_module_monitor module_monitor_68;
    nodf_module_intf module_intf_69(clock,reset);
    assign module_intf_69.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.call_ln212_write_p4_fu_153.ap_start;
    assign module_intf_69.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.call_ln212_write_p4_fu_153.ap_ready;
    assign module_intf_69.ap_done = 1'b0;
    assign module_intf_69.ap_continue = 1'b0;
    assign module_intf_69.finish = finish;
    csv_file_dump mstatus_csv_dumper_69;
    nodf_module_monitor module_monitor_69;
    nodf_module_intf module_intf_70(clock,reset);
    assign module_intf_70.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_start;
    assign module_intf_70.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_ready;
    assign module_intf_70.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_done;
    assign module_intf_70.ap_continue = 1'b1;
    assign module_intf_70.finish = finish;
    csv_file_dump mstatus_csv_dumper_70;
    nodf_module_monitor module_monitor_70;
    nodf_module_intf module_intf_71(clock,reset);
    assign module_intf_71.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.grp_read_p1_fu_164.ap_start;
    assign module_intf_71.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.grp_read_p1_fu_164.ap_ready;
    assign module_intf_71.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.grp_read_p1_fu_164.ap_done;
    assign module_intf_71.ap_continue = 1'b1;
    assign module_intf_71.finish = finish;
    csv_file_dump mstatus_csv_dumper_71;
    nodf_module_monitor module_monitor_71;
    nodf_module_intf module_intf_72(clock,reset);
    assign module_intf_72.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.grp_read_p2_fu_171.ap_start;
    assign module_intf_72.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.grp_read_p2_fu_171.ap_ready;
    assign module_intf_72.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.grp_read_p2_fu_171.ap_done;
    assign module_intf_72.ap_continue = 1'b1;
    assign module_intf_72.finish = finish;
    csv_file_dump mstatus_csv_dumper_72;
    nodf_module_monitor module_monitor_72;
    nodf_module_intf module_intf_73(clock,reset);
    assign module_intf_73.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.call_ln221_write_p3_fu_187.ap_start;
    assign module_intf_73.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.call_ln221_write_p3_fu_187.ap_ready;
    assign module_intf_73.ap_done = 1'b0;
    assign module_intf_73.ap_continue = 1'b0;
    assign module_intf_73.finish = finish;
    csv_file_dump mstatus_csv_dumper_73;
    nodf_module_monitor module_monitor_73;
    nodf_module_intf module_intf_74(clock,reset);
    assign module_intf_74.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_start;
    assign module_intf_74.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_ready;
    assign module_intf_74.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_done;
    assign module_intf_74.ap_continue = 1'b1;
    assign module_intf_74.finish = finish;
    csv_file_dump mstatus_csv_dumper_74;
    nodf_module_monitor module_monitor_74;
    nodf_module_intf module_intf_75(clock,reset);
    assign module_intf_75.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.grp_read_p1_fu_137.ap_start;
    assign module_intf_75.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.grp_read_p1_fu_137.ap_ready;
    assign module_intf_75.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.grp_read_p1_fu_137.ap_done;
    assign module_intf_75.ap_continue = 1'b1;
    assign module_intf_75.finish = finish;
    csv_file_dump mstatus_csv_dumper_75;
    nodf_module_monitor module_monitor_75;
    nodf_module_intf module_intf_76(clock,reset);
    assign module_intf_76.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.call_ln173_write_p3_fu_153.ap_start;
    assign module_intf_76.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.call_ln173_write_p3_fu_153.ap_ready;
    assign module_intf_76.ap_done = 1'b0;
    assign module_intf_76.ap_continue = 1'b0;
    assign module_intf_76.finish = finish;
    csv_file_dump mstatus_csv_dumper_76;
    nodf_module_monitor module_monitor_76;
    nodf_module_intf module_intf_77(clock,reset);
    assign module_intf_77.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_start;
    assign module_intf_77.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_ready;
    assign module_intf_77.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_done;
    assign module_intf_77.ap_continue = 1'b1;
    assign module_intf_77.finish = finish;
    csv_file_dump mstatus_csv_dumper_77;
    nodf_module_monitor module_monitor_77;
    nodf_module_intf module_intf_78(clock,reset);
    assign module_intf_78.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.grp_read_p1_fu_162.ap_start;
    assign module_intf_78.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.grp_read_p1_fu_162.ap_ready;
    assign module_intf_78.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.grp_read_p1_fu_162.ap_done;
    assign module_intf_78.ap_continue = 1'b1;
    assign module_intf_78.finish = finish;
    csv_file_dump mstatus_csv_dumper_78;
    nodf_module_monitor module_monitor_78;
    nodf_module_intf module_intf_79(clock,reset);
    assign module_intf_79.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.grp_read_p2_fu_169.ap_start;
    assign module_intf_79.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.grp_read_p2_fu_169.ap_ready;
    assign module_intf_79.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.grp_read_p2_fu_169.ap_done;
    assign module_intf_79.ap_continue = 1'b1;
    assign module_intf_79.finish = finish;
    csv_file_dump mstatus_csv_dumper_79;
    nodf_module_monitor module_monitor_79;
    nodf_module_intf module_intf_80(clock,reset);
    assign module_intf_80.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.call_ln182_write_p3_fu_185.ap_start;
    assign module_intf_80.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.call_ln182_write_p3_fu_185.ap_ready;
    assign module_intf_80.ap_done = 1'b0;
    assign module_intf_80.ap_continue = 1'b0;
    assign module_intf_80.finish = finish;
    csv_file_dump mstatus_csv_dumper_80;
    nodf_module_monitor module_monitor_80;
    nodf_module_intf module_intf_81(clock,reset);
    assign module_intf_81.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_start;
    assign module_intf_81.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_ready;
    assign module_intf_81.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_done;
    assign module_intf_81.ap_continue = 1'b1;
    assign module_intf_81.finish = finish;
    csv_file_dump mstatus_csv_dumper_81;
    nodf_module_monitor module_monitor_81;
    nodf_module_intf module_intf_82(clock,reset);
    assign module_intf_82.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.grp_read_intt_fu_137.ap_start;
    assign module_intf_82.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.grp_read_intt_fu_137.ap_ready;
    assign module_intf_82.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.grp_read_intt_fu_137.ap_done;
    assign module_intf_82.ap_continue = 1'b1;
    assign module_intf_82.finish = finish;
    csv_file_dump mstatus_csv_dumper_82;
    nodf_module_monitor module_monitor_82;
    nodf_module_intf module_intf_83(clock,reset);
    assign module_intf_83.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.call_ln350_write_p3_fu_153.ap_start;
    assign module_intf_83.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.call_ln350_write_p3_fu_153.ap_ready;
    assign module_intf_83.ap_done = 1'b0;
    assign module_intf_83.ap_continue = 1'b0;
    assign module_intf_83.finish = finish;
    csv_file_dump mstatus_csv_dumper_83;
    nodf_module_monitor module_monitor_83;
    nodf_module_intf module_intf_84(clock,reset);
    assign module_intf_84.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_start;
    assign module_intf_84.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_ready;
    assign module_intf_84.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_done;
    assign module_intf_84.ap_continue = 1'b1;
    assign module_intf_84.finish = finish;
    csv_file_dump mstatus_csv_dumper_84;
    nodf_module_monitor module_monitor_84;
    nodf_module_intf module_intf_85(clock,reset);
    assign module_intf_85.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.grp_read_p1_fu_151.ap_start;
    assign module_intf_85.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.grp_read_p1_fu_151.ap_ready;
    assign module_intf_85.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.grp_read_p1_fu_151.ap_done;
    assign module_intf_85.ap_continue = 1'b1;
    assign module_intf_85.finish = finish;
    csv_file_dump mstatus_csv_dumper_85;
    nodf_module_monitor module_monitor_85;
    nodf_module_intf module_intf_86(clock,reset);
    assign module_intf_86.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.call_ln358_write_p3_fu_167.ap_start;
    assign module_intf_86.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.call_ln358_write_p3_fu_167.ap_ready;
    assign module_intf_86.ap_done = 1'b0;
    assign module_intf_86.ap_continue = 1'b0;
    assign module_intf_86.finish = finish;
    csv_file_dump mstatus_csv_dumper_86;
    nodf_module_monitor module_monitor_86;
    nodf_module_intf module_intf_87(clock,reset);
    assign module_intf_87.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.call_ln359_write_p4_fu_175.ap_start;
    assign module_intf_87.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.call_ln359_write_p4_fu_175.ap_ready;
    assign module_intf_87.ap_done = 1'b0;
    assign module_intf_87.ap_continue = 1'b0;
    assign module_intf_87.finish = finish;
    csv_file_dump mstatus_csv_dumper_87;
    nodf_module_monitor module_monitor_87;
    nodf_module_intf module_intf_88(clock,reset);
    assign module_intf_88.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_start;
    assign module_intf_88.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_ready;
    assign module_intf_88.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_done;
    assign module_intf_88.ap_continue = 1'b1;
    assign module_intf_88.finish = finish;
    csv_file_dump mstatus_csv_dumper_88;
    nodf_module_monitor module_monitor_88;
    nodf_module_intf module_intf_89(clock,reset);
    assign module_intf_89.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.grp_read_p1_fu_137.ap_start;
    assign module_intf_89.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.grp_read_p1_fu_137.ap_ready;
    assign module_intf_89.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.grp_read_p1_fu_137.ap_done;
    assign module_intf_89.ap_continue = 1'b1;
    assign module_intf_89.finish = finish;
    csv_file_dump mstatus_csv_dumper_89;
    nodf_module_monitor module_monitor_89;
    nodf_module_intf module_intf_90(clock,reset);
    assign module_intf_90.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.call_ln368_write_p3_fu_153.ap_start;
    assign module_intf_90.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.call_ln368_write_p3_fu_153.ap_ready;
    assign module_intf_90.ap_done = 1'b0;
    assign module_intf_90.ap_continue = 1'b0;
    assign module_intf_90.finish = finish;
    csv_file_dump mstatus_csv_dumper_90;
    nodf_module_monitor module_monitor_90;
    nodf_module_intf module_intf_91(clock,reset);
    assign module_intf_91.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_start;
    assign module_intf_91.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_ready;
    assign module_intf_91.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_done;
    assign module_intf_91.ap_continue = 1'b1;
    assign module_intf_91.finish = finish;
    csv_file_dump mstatus_csv_dumper_91;
    nodf_module_monitor module_monitor_91;
    nodf_module_intf module_intf_92(clock,reset);
    assign module_intf_92.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.grp_read_p1_fu_137.ap_start;
    assign module_intf_92.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.grp_read_p1_fu_137.ap_ready;
    assign module_intf_92.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.grp_read_p1_fu_137.ap_done;
    assign module_intf_92.ap_continue = 1'b1;
    assign module_intf_92.finish = finish;
    csv_file_dump mstatus_csv_dumper_92;
    nodf_module_monitor module_monitor_92;
    nodf_module_intf module_intf_93(clock,reset);
    assign module_intf_93.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.call_ln377_write_p4_fu_153.ap_start;
    assign module_intf_93.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.call_ln377_write_p4_fu_153.ap_ready;
    assign module_intf_93.ap_done = 1'b0;
    assign module_intf_93.ap_continue = 1'b0;
    assign module_intf_93.finish = finish;
    csv_file_dump mstatus_csv_dumper_93;
    nodf_module_monitor module_monitor_93;
    nodf_module_intf module_intf_94(clock,reset);
    assign module_intf_94.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_start;
    assign module_intf_94.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_ready;
    assign module_intf_94.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_done;
    assign module_intf_94.ap_continue = 1'b1;
    assign module_intf_94.finish = finish;
    csv_file_dump mstatus_csv_dumper_94;
    nodf_module_monitor module_monitor_94;
    nodf_module_intf module_intf_95(clock,reset);
    assign module_intf_95.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.grp_read_p1_fu_118.ap_start;
    assign module_intf_95.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.grp_read_p1_fu_118.ap_ready;
    assign module_intf_95.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.grp_read_p1_fu_118.ap_done;
    assign module_intf_95.ap_continue = 1'b1;
    assign module_intf_95.finish = finish;
    csv_file_dump mstatus_csv_dumper_95;
    nodf_module_monitor module_monitor_95;
    nodf_module_intf module_intf_96(clock,reset);
    assign module_intf_96.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.grp_read_p2_fu_125.ap_start;
    assign module_intf_96.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.grp_read_p2_fu_125.ap_ready;
    assign module_intf_96.ap_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.grp_read_p2_fu_125.ap_done;
    assign module_intf_96.ap_continue = 1'b1;
    assign module_intf_96.finish = finish;
    csv_file_dump mstatus_csv_dumper_96;
    nodf_module_monitor module_monitor_96;
    nodf_module_intf module_intf_97(clock,reset);
    assign module_intf_97.ap_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.call_ln386_write_p3_fu_141.ap_start;
    assign module_intf_97.ap_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.call_ln386_write_p3_fu_141.ap_ready;
    assign module_intf_97.ap_done = 1'b0;
    assign module_intf_97.ap_continue = 1'b0;
    assign module_intf_97.finish = finish;
    csv_file_dump mstatus_csv_dumper_97;
    nodf_module_monitor module_monitor_97;
    nodf_module_intf module_intf_98(clock,reset);
    assign module_intf_98.ap_start = 1'b0;
    assign module_intf_98.ap_ready = 1'b0;
    assign module_intf_98.ap_done = 1'b0;
    assign module_intf_98.ap_continue = 1'b0;
    assign module_intf_98.finish = finish;
    csv_file_dump mstatus_csv_dumper_98;
    nodf_module_monitor module_monitor_98;
    nodf_module_intf module_intf_99(clock,reset);
    assign module_intf_99.ap_start = 1'b0;
    assign module_intf_99.ap_ready = 1'b0;
    assign module_intf_99.ap_done = 1'b0;
    assign module_intf_99.ap_continue = 1'b0;
    assign module_intf_99.finish = finish;
    csv_file_dump mstatus_csv_dumper_99;
    nodf_module_monitor module_monitor_99;
    nodf_module_intf module_intf_100(clock,reset);
    assign module_intf_100.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_40_1_fu_562.ap_start;
    assign module_intf_100.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_40_1_fu_562.ap_ready;
    assign module_intf_100.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_40_1_fu_562.ap_done;
    assign module_intf_100.ap_continue = 1'b1;
    assign module_intf_100.finish = finish;
    csv_file_dump mstatus_csv_dumper_100;
    nodf_module_monitor module_monitor_100;
    nodf_module_intf module_intf_101(clock,reset);
    assign module_intf_101.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_41_2_fu_567.ap_start;
    assign module_intf_101.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_41_2_fu_567.ap_ready;
    assign module_intf_101.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_41_2_fu_567.ap_done;
    assign module_intf_101.ap_continue = 1'b1;
    assign module_intf_101.finish = finish;
    csv_file_dump mstatus_csv_dumper_101;
    nodf_module_monitor module_monitor_101;
    nodf_module_intf module_intf_102(clock,reset);
    assign module_intf_102.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_1_fu_572.ap_start;
    assign module_intf_102.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_1_fu_572.ap_ready;
    assign module_intf_102.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_1_fu_572.ap_done;
    assign module_intf_102.ap_continue = 1'b1;
    assign module_intf_102.finish = finish;
    csv_file_dump mstatus_csv_dumper_102;
    nodf_module_monitor module_monitor_102;
    nodf_module_intf module_intf_103(clock,reset);
    assign module_intf_103.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_start;
    assign module_intf_103.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_ready;
    assign module_intf_103.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_done;
    assign module_intf_103.ap_continue = 1'b1;
    assign module_intf_103.finish = finish;
    csv_file_dump mstatus_csv_dumper_103;
    nodf_module_monitor module_monitor_103;
    nodf_module_intf module_intf_104(clock,reset);
    assign module_intf_104.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_start;
    assign module_intf_104.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ready;
    assign module_intf_104.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_done;
    assign module_intf_104.ap_continue = 1'b1;
    assign module_intf_104.finish = finish;
    csv_file_dump mstatus_csv_dumper_104;
    nodf_module_monitor module_monitor_104;
    nodf_module_intf module_intf_105(clock,reset);
    assign module_intf_105.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_start;
    assign module_intf_105.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ready;
    assign module_intf_105.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_done;
    assign module_intf_105.ap_continue = 1'b1;
    assign module_intf_105.finish = finish;
    csv_file_dump mstatus_csv_dumper_105;
    nodf_module_monitor module_monitor_105;
    nodf_module_intf module_intf_106(clock,reset);
    assign module_intf_106.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_start;
    assign module_intf_106.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ready;
    assign module_intf_106.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_done;
    assign module_intf_106.ap_continue = 1'b1;
    assign module_intf_106.finish = finish;
    csv_file_dump mstatus_csv_dumper_106;
    nodf_module_monitor module_monitor_106;
    nodf_module_intf module_intf_107(clock,reset);
    assign module_intf_107.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_start;
    assign module_intf_107.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_ready;
    assign module_intf_107.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_done;
    assign module_intf_107.ap_continue = 1'b1;
    assign module_intf_107.finish = finish;
    csv_file_dump mstatus_csv_dumper_107;
    nodf_module_monitor module_monitor_107;
    nodf_module_intf module_intf_108(clock,reset);
    assign module_intf_108.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_383_6_fu_172.ap_start;
    assign module_intf_108.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_383_6_fu_172.ap_ready;
    assign module_intf_108.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_383_6_fu_172.ap_done;
    assign module_intf_108.ap_continue = 1'b1;
    assign module_intf_108.finish = finish;
    csv_file_dump mstatus_csv_dumper_108;
    nodf_module_monitor module_monitor_108;
    nodf_module_intf module_intf_109(clock,reset);
    assign module_intf_109.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_start;
    assign module_intf_109.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ready;
    assign module_intf_109.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_done;
    assign module_intf_109.ap_continue = 1'b1;
    assign module_intf_109.finish = finish;
    csv_file_dump mstatus_csv_dumper_109;
    nodf_module_monitor module_monitor_109;
    nodf_module_intf module_intf_110(clock,reset);
    assign module_intf_110.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_start;
    assign module_intf_110.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ready;
    assign module_intf_110.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_done;
    assign module_intf_110.ap_continue = 1'b1;
    assign module_intf_110.finish = finish;
    csv_file_dump mstatus_csv_dumper_110;
    nodf_module_monitor module_monitor_110;
    nodf_module_intf module_intf_111(clock,reset);
    assign module_intf_111.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_start;
    assign module_intf_111.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_ready;
    assign module_intf_111.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_done;
    assign module_intf_111.ap_continue = 1'b1;
    assign module_intf_111.finish = finish;
    csv_file_dump mstatus_csv_dumper_111;
    nodf_module_monitor module_monitor_111;
    nodf_module_intf module_intf_112(clock,reset);
    assign module_intf_112.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_start;
    assign module_intf_112.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_ready;
    assign module_intf_112.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_done;
    assign module_intf_112.ap_continue = 1'b1;
    assign module_intf_112.finish = finish;
    csv_file_dump mstatus_csv_dumper_112;
    nodf_module_monitor module_monitor_112;
    nodf_module_intf module_intf_113(clock,reset);
    assign module_intf_113.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_start;
    assign module_intf_113.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_ready;
    assign module_intf_113.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_done;
    assign module_intf_113.ap_continue = 1'b1;
    assign module_intf_113.finish = finish;
    csv_file_dump mstatus_csv_dumper_113;
    nodf_module_monitor module_monitor_113;
    nodf_module_intf module_intf_114(clock,reset);
    assign module_intf_114.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_start;
    assign module_intf_114.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_ready;
    assign module_intf_114.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_done;
    assign module_intf_114.ap_continue = 1'b1;
    assign module_intf_114.finish = finish;
    csv_file_dump mstatus_csv_dumper_114;
    nodf_module_monitor module_monitor_114;
    nodf_module_intf module_intf_115(clock,reset);
    assign module_intf_115.ap_start = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_start;
    assign module_intf_115.ap_ready = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_ready;
    assign module_intf_115.ap_done = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_done;
    assign module_intf_115.ap_continue = 1'b1;
    assign module_intf_115.finish = finish;
    csv_file_dump mstatus_csv_dumper_115;
    nodf_module_monitor module_monitor_115;
    nodf_module_intf module_intf_116(clock,reset);
    assign module_intf_116.ap_start = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_start;
    assign module_intf_116.ap_ready = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_ready;
    assign module_intf_116.ap_done = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_done;
    assign module_intf_116.ap_continue = 1'b1;
    assign module_intf_116.finish = finish;
    csv_file_dump mstatus_csv_dumper_116;
    nodf_module_monitor module_monitor_116;
    nodf_module_intf module_intf_117(clock,reset);
    assign module_intf_117.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_16_fu_635.ap_start;
    assign module_intf_117.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_16_fu_635.ap_ready;
    assign module_intf_117.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_16_fu_635.ap_done;
    assign module_intf_117.ap_continue = 1'b1;
    assign module_intf_117.finish = finish;
    csv_file_dump mstatus_csv_dumper_117;
    nodf_module_monitor module_monitor_117;
    nodf_module_intf module_intf_118(clock,reset);
    assign module_intf_118.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_start;
    assign module_intf_118.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ready;
    assign module_intf_118.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_done;
    assign module_intf_118.ap_continue = 1'b1;
    assign module_intf_118.finish = finish;
    csv_file_dump mstatus_csv_dumper_118;
    nodf_module_monitor module_monitor_118;
    nodf_module_intf module_intf_119(clock,reset);
    assign module_intf_119.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_start;
    assign module_intf_119.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ready;
    assign module_intf_119.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_done;
    assign module_intf_119.ap_continue = 1'b1;
    assign module_intf_119.finish = finish;
    csv_file_dump mstatus_csv_dumper_119;
    nodf_module_monitor module_monitor_119;
    nodf_module_intf module_intf_120(clock,reset);
    assign module_intf_120.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_start;
    assign module_intf_120.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ready;
    assign module_intf_120.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_done;
    assign module_intf_120.ap_continue = 1'b1;
    assign module_intf_120.finish = finish;
    csv_file_dump mstatus_csv_dumper_120;
    nodf_module_monitor module_monitor_120;
    nodf_module_intf module_intf_121(clock,reset);
    assign module_intf_121.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_start;
    assign module_intf_121.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ready;
    assign module_intf_121.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_done;
    assign module_intf_121.ap_continue = 1'b1;
    assign module_intf_121.finish = finish;
    csv_file_dump mstatus_csv_dumper_121;
    nodf_module_monitor module_monitor_121;
    nodf_module_intf module_intf_122(clock,reset);
    assign module_intf_122.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_start;
    assign module_intf_122.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_ready;
    assign module_intf_122.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_done;
    assign module_intf_122.ap_continue = 1'b1;
    assign module_intf_122.finish = finish;
    csv_file_dump mstatus_csv_dumper_122;
    nodf_module_monitor module_monitor_122;
    nodf_module_intf module_intf_123(clock,reset);
    assign module_intf_123.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_start;
    assign module_intf_123.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ready;
    assign module_intf_123.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_done;
    assign module_intf_123.ap_continue = 1'b1;
    assign module_intf_123.finish = finish;
    csv_file_dump mstatus_csv_dumper_123;
    nodf_module_monitor module_monitor_123;
    nodf_module_intf module_intf_124(clock,reset);
    assign module_intf_124.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_start;
    assign module_intf_124.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ready;
    assign module_intf_124.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_done;
    assign module_intf_124.ap_continue = 1'b1;
    assign module_intf_124.finish = finish;
    csv_file_dump mstatus_csv_dumper_124;
    nodf_module_monitor module_monitor_124;
    nodf_module_intf module_intf_125(clock,reset);
    assign module_intf_125.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_383_6_fu_293.ap_start;
    assign module_intf_125.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_383_6_fu_293.ap_ready;
    assign module_intf_125.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_383_6_fu_293.ap_done;
    assign module_intf_125.ap_continue = 1'b1;
    assign module_intf_125.finish = finish;
    csv_file_dump mstatus_csv_dumper_125;
    nodf_module_monitor module_monitor_125;
    nodf_module_intf module_intf_126(clock,reset);
    assign module_intf_126.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_385_7_fu_298.ap_start;
    assign module_intf_126.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_385_7_fu_298.ap_ready;
    assign module_intf_126.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_385_7_fu_298.ap_done;
    assign module_intf_126.ap_continue = 1'b1;
    assign module_intf_126.finish = finish;
    csv_file_dump mstatus_csv_dumper_126;
    nodf_module_monitor module_monitor_126;
    nodf_module_intf module_intf_127(clock,reset);
    assign module_intf_127.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_start;
    assign module_intf_127.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ready;
    assign module_intf_127.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_done;
    assign module_intf_127.ap_continue = 1'b1;
    assign module_intf_127.finish = finish;
    csv_file_dump mstatus_csv_dumper_127;
    nodf_module_monitor module_monitor_127;
    nodf_module_intf module_intf_128(clock,reset);
    assign module_intf_128.ap_start = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_start;
    assign module_intf_128.ap_ready = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_ready;
    assign module_intf_128.ap_done = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_done;
    assign module_intf_128.ap_continue = 1'b1;
    assign module_intf_128.finish = finish;
    csv_file_dump mstatus_csv_dumper_128;
    nodf_module_monitor module_monitor_128;
    nodf_module_intf module_intf_129(clock,reset);
    assign module_intf_129.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_start;
    assign module_intf_129.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_ready;
    assign module_intf_129.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_done;
    assign module_intf_129.ap_continue = 1'b1;
    assign module_intf_129.finish = finish;
    csv_file_dump mstatus_csv_dumper_129;
    nodf_module_monitor module_monitor_129;
    nodf_module_intf module_intf_130(clock,reset);
    assign module_intf_130.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_start;
    assign module_intf_130.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_ready;
    assign module_intf_130.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_done;
    assign module_intf_130.ap_continue = 1'b1;
    assign module_intf_130.finish = finish;
    csv_file_dump mstatus_csv_dumper_130;
    nodf_module_monitor module_monitor_130;
    nodf_module_intf module_intf_131(clock,reset);
    assign module_intf_131.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_start;
    assign module_intf_131.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_ready;
    assign module_intf_131.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_done;
    assign module_intf_131.ap_continue = 1'b1;
    assign module_intf_131.finish = finish;
    csv_file_dump mstatus_csv_dumper_131;
    nodf_module_monitor module_monitor_131;
    nodf_module_intf module_intf_132(clock,reset);
    assign module_intf_132.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_start;
    assign module_intf_132.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ready;
    assign module_intf_132.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_done;
    assign module_intf_132.ap_continue = 1'b1;
    assign module_intf_132.finish = finish;
    csv_file_dump mstatus_csv_dumper_132;
    nodf_module_monitor module_monitor_132;
    nodf_module_intf module_intf_133(clock,reset);
    assign module_intf_133.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_start;
    assign module_intf_133.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ready;
    assign module_intf_133.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_done;
    assign module_intf_133.ap_continue = 1'b1;
    assign module_intf_133.finish = finish;
    csv_file_dump mstatus_csv_dumper_133;
    nodf_module_monitor module_monitor_133;
    nodf_module_intf module_intf_134(clock,reset);
    assign module_intf_134.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_start;
    assign module_intf_134.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ready;
    assign module_intf_134.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_done;
    assign module_intf_134.ap_continue = 1'b1;
    assign module_intf_134.finish = finish;
    csv_file_dump mstatus_csv_dumper_134;
    nodf_module_monitor module_monitor_134;
    nodf_module_intf module_intf_135(clock,reset);
    assign module_intf_135.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_start;
    assign module_intf_135.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ready;
    assign module_intf_135.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_done;
    assign module_intf_135.ap_continue = 1'b1;
    assign module_intf_135.finish = finish;
    csv_file_dump mstatus_csv_dumper_135;
    nodf_module_monitor module_monitor_135;
    nodf_module_intf module_intf_136(clock,reset);
    assign module_intf_136.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_start;
    assign module_intf_136.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_ready;
    assign module_intf_136.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_done;
    assign module_intf_136.ap_continue = 1'b1;
    assign module_intf_136.finish = finish;
    csv_file_dump mstatus_csv_dumper_136;
    nodf_module_monitor module_monitor_136;
    nodf_module_intf module_intf_137(clock,reset);
    assign module_intf_137.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_383_6_fu_172.ap_start;
    assign module_intf_137.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_383_6_fu_172.ap_ready;
    assign module_intf_137.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_383_6_fu_172.ap_done;
    assign module_intf_137.ap_continue = 1'b1;
    assign module_intf_137.finish = finish;
    csv_file_dump mstatus_csv_dumper_137;
    nodf_module_monitor module_monitor_137;
    nodf_module_intf module_intf_138(clock,reset);
    assign module_intf_138.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_start;
    assign module_intf_138.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ready;
    assign module_intf_138.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_done;
    assign module_intf_138.ap_continue = 1'b1;
    assign module_intf_138.finish = finish;
    csv_file_dump mstatus_csv_dumper_138;
    nodf_module_monitor module_monitor_138;
    nodf_module_intf module_intf_139(clock,reset);
    assign module_intf_139.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_start;
    assign module_intf_139.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ready;
    assign module_intf_139.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_done;
    assign module_intf_139.ap_continue = 1'b1;
    assign module_intf_139.finish = finish;
    csv_file_dump mstatus_csv_dumper_139;
    nodf_module_monitor module_monitor_139;
    nodf_module_intf module_intf_140(clock,reset);
    assign module_intf_140.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_start;
    assign module_intf_140.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ready;
    assign module_intf_140.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_done;
    assign module_intf_140.ap_continue = 1'b1;
    assign module_intf_140.finish = finish;
    csv_file_dump mstatus_csv_dumper_140;
    nodf_module_monitor module_monitor_140;
    nodf_module_intf module_intf_141(clock,reset);
    assign module_intf_141.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_start;
    assign module_intf_141.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ready;
    assign module_intf_141.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_done;
    assign module_intf_141.ap_continue = 1'b1;
    assign module_intf_141.finish = finish;
    csv_file_dump mstatus_csv_dumper_141;
    nodf_module_monitor module_monitor_141;
    nodf_module_intf module_intf_142(clock,reset);
    assign module_intf_142.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_start;
    assign module_intf_142.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ready;
    assign module_intf_142.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_done;
    assign module_intf_142.ap_continue = 1'b1;
    assign module_intf_142.finish = finish;
    csv_file_dump mstatus_csv_dumper_142;
    nodf_module_monitor module_monitor_142;
    nodf_module_intf module_intf_143(clock,reset);
    assign module_intf_143.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_start;
    assign module_intf_143.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ready;
    assign module_intf_143.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_done;
    assign module_intf_143.ap_continue = 1'b1;
    assign module_intf_143.finish = finish;
    csv_file_dump mstatus_csv_dumper_143;
    nodf_module_monitor module_monitor_143;
    nodf_module_intf module_intf_144(clock,reset);
    assign module_intf_144.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_start;
    assign module_intf_144.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_ready;
    assign module_intf_144.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_done;
    assign module_intf_144.ap_continue = 1'b1;
    assign module_intf_144.finish = finish;
    csv_file_dump mstatus_csv_dumper_144;
    nodf_module_monitor module_monitor_144;
    nodf_module_intf module_intf_145(clock,reset);
    assign module_intf_145.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_start;
    assign module_intf_145.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ready;
    assign module_intf_145.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_done;
    assign module_intf_145.ap_continue = 1'b1;
    assign module_intf_145.finish = finish;
    csv_file_dump mstatus_csv_dumper_145;
    nodf_module_monitor module_monitor_145;
    nodf_module_intf module_intf_146(clock,reset);
    assign module_intf_146.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_start;
    assign module_intf_146.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ready;
    assign module_intf_146.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_done;
    assign module_intf_146.ap_continue = 1'b1;
    assign module_intf_146.finish = finish;
    csv_file_dump mstatus_csv_dumper_146;
    nodf_module_monitor module_monitor_146;
    nodf_module_intf module_intf_147(clock,reset);
    assign module_intf_147.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_383_6_fu_293.ap_start;
    assign module_intf_147.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_383_6_fu_293.ap_ready;
    assign module_intf_147.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_383_6_fu_293.ap_done;
    assign module_intf_147.ap_continue = 1'b1;
    assign module_intf_147.finish = finish;
    csv_file_dump mstatus_csv_dumper_147;
    nodf_module_monitor module_monitor_147;
    nodf_module_intf module_intf_148(clock,reset);
    assign module_intf_148.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_385_7_fu_298.ap_start;
    assign module_intf_148.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_385_7_fu_298.ap_ready;
    assign module_intf_148.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_385_7_fu_298.ap_done;
    assign module_intf_148.ap_continue = 1'b1;
    assign module_intf_148.finish = finish;
    csv_file_dump mstatus_csv_dumper_148;
    nodf_module_monitor module_monitor_148;
    nodf_module_intf module_intf_149(clock,reset);
    assign module_intf_149.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_start;
    assign module_intf_149.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ready;
    assign module_intf_149.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_done;
    assign module_intf_149.ap_continue = 1'b1;
    assign module_intf_149.finish = finish;
    csv_file_dump mstatus_csv_dumper_149;
    nodf_module_monitor module_monitor_149;
    nodf_module_intf module_intf_150(clock,reset);
    assign module_intf_150.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_start;
    assign module_intf_150.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_ready;
    assign module_intf_150.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_done;
    assign module_intf_150.ap_continue = 1'b1;
    assign module_intf_150.finish = finish;
    csv_file_dump mstatus_csv_dumper_150;
    nodf_module_monitor module_monitor_150;
    nodf_module_intf module_intf_151(clock,reset);
    assign module_intf_151.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_start;
    assign module_intf_151.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_ready;
    assign module_intf_151.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_done;
    assign module_intf_151.ap_continue = 1'b1;
    assign module_intf_151.finish = finish;
    csv_file_dump mstatus_csv_dumper_151;
    nodf_module_monitor module_monitor_151;
    nodf_module_intf module_intf_152(clock,reset);
    assign module_intf_152.ap_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_start;
    assign module_intf_152.ap_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_ready;
    assign module_intf_152.ap_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_done;
    assign module_intf_152.ap_continue = 1'b1;
    assign module_intf_152.finish = finish;
    csv_file_dump mstatus_csv_dumper_152;
    nodf_module_monitor module_monitor_152;
    nodf_module_intf module_intf_153(clock,reset);
    assign module_intf_153.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_start;
    assign module_intf_153.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_ready;
    assign module_intf_153.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_done;
    assign module_intf_153.ap_continue = 1'b1;
    assign module_intf_153.finish = finish;
    csv_file_dump mstatus_csv_dumper_153;
    nodf_module_monitor module_monitor_153;
    nodf_module_intf module_intf_154(clock,reset);
    assign module_intf_154.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_start;
    assign module_intf_154.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_ready;
    assign module_intf_154.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_done;
    assign module_intf_154.ap_continue = 1'b1;
    assign module_intf_154.finish = finish;
    csv_file_dump mstatus_csv_dumper_154;
    nodf_module_monitor module_monitor_154;
    nodf_module_intf module_intf_155(clock,reset);
    assign module_intf_155.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_start;
    assign module_intf_155.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_ready;
    assign module_intf_155.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_done;
    assign module_intf_155.ap_continue = 1'b1;
    assign module_intf_155.finish = finish;
    csv_file_dump mstatus_csv_dumper_155;
    nodf_module_monitor module_monitor_155;
    nodf_module_intf module_intf_156(clock,reset);
    assign module_intf_156.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_110_fu_714.ap_start;
    assign module_intf_156.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_110_fu_714.ap_ready;
    assign module_intf_156.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_321_110_fu_714.ap_done;
    assign module_intf_156.ap_continue = 1'b1;
    assign module_intf_156.finish = finish;
    csv_file_dump mstatus_csv_dumper_156;
    nodf_module_monitor module_monitor_156;
    nodf_module_intf module_intf_157(clock,reset);
    assign module_intf_157.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_start;
    assign module_intf_157.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_ready;
    assign module_intf_157.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_done;
    assign module_intf_157.ap_continue = 1'b1;
    assign module_intf_157.finish = finish;
    csv_file_dump mstatus_csv_dumper_157;
    nodf_module_monitor module_monitor_157;
    nodf_module_intf module_intf_158(clock,reset);
    assign module_intf_158.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_start;
    assign module_intf_158.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_ready;
    assign module_intf_158.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_done;
    assign module_intf_158.ap_continue = 1'b1;
    assign module_intf_158.finish = finish;
    csv_file_dump mstatus_csv_dumper_158;
    nodf_module_monitor module_monitor_158;
    nodf_module_intf module_intf_159(clock,reset);
    assign module_intf_159.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_start;
    assign module_intf_159.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_ready;
    assign module_intf_159.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_done;
    assign module_intf_159.ap_continue = 1'b1;
    assign module_intf_159.finish = finish;
    csv_file_dump mstatus_csv_dumper_159;
    nodf_module_monitor module_monitor_159;
    nodf_module_intf module_intf_160(clock,reset);
    assign module_intf_160.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_start;
    assign module_intf_160.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_ready;
    assign module_intf_160.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_done;
    assign module_intf_160.ap_continue = 1'b1;
    assign module_intf_160.finish = finish;
    csv_file_dump mstatus_csv_dumper_160;
    nodf_module_monitor module_monitor_160;
    nodf_module_intf module_intf_161(clock,reset);
    assign module_intf_161.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_start;
    assign module_intf_161.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_ready;
    assign module_intf_161.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_done;
    assign module_intf_161.ap_continue = 1'b1;
    assign module_intf_161.finish = finish;
    csv_file_dump mstatus_csv_dumper_161;
    nodf_module_monitor module_monitor_161;
    nodf_module_intf module_intf_162(clock,reset);
    assign module_intf_162.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_605_2_fu_87.ap_start;
    assign module_intf_162.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_605_2_fu_87.ap_ready;
    assign module_intf_162.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_605_2_fu_87.ap_done;
    assign module_intf_162.ap_continue = 1'b1;
    assign module_intf_162.finish = finish;
    csv_file_dump mstatus_csv_dumper_162;
    nodf_module_monitor module_monitor_162;
    nodf_module_intf module_intf_163(clock,reset);
    assign module_intf_163.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_start;
    assign module_intf_163.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_ready;
    assign module_intf_163.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_done;
    assign module_intf_163.ap_continue = 1'b1;
    assign module_intf_163.finish = finish;
    csv_file_dump mstatus_csv_dumper_163;
    nodf_module_monitor module_monitor_163;
    nodf_module_intf module_intf_164(clock,reset);
    assign module_intf_164.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_start;
    assign module_intf_164.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_ready;
    assign module_intf_164.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_done;
    assign module_intf_164.ap_continue = 1'b1;
    assign module_intf_164.finish = finish;
    csv_file_dump mstatus_csv_dumper_164;
    nodf_module_monitor module_monitor_164;
    nodf_module_intf module_intf_165(clock,reset);
    assign module_intf_165.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_start;
    assign module_intf_165.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_ready;
    assign module_intf_165.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_done;
    assign module_intf_165.ap_continue = 1'b1;
    assign module_intf_165.finish = finish;
    csv_file_dump mstatus_csv_dumper_165;
    nodf_module_monitor module_monitor_165;
    nodf_module_intf module_intf_166(clock,reset);
    assign module_intf_166.ap_start = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_start;
    assign module_intf_166.ap_ready = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_ready;
    assign module_intf_166.ap_done = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_done;
    assign module_intf_166.ap_continue = 1'b1;
    assign module_intf_166.finish = finish;
    csv_file_dump mstatus_csv_dumper_166;
    nodf_module_monitor module_monitor_166;
    nodf_module_intf module_intf_167(clock,reset);
    assign module_intf_167.ap_start = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_start;
    assign module_intf_167.ap_ready = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_ready;
    assign module_intf_167.ap_done = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_done;
    assign module_intf_167.ap_continue = 1'b1;
    assign module_intf_167.finish = finish;
    csv_file_dump mstatus_csv_dumper_167;
    nodf_module_monitor module_monitor_167;
    nodf_module_intf module_intf_168(clock,reset);
    assign module_intf_168.ap_start = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_start;
    assign module_intf_168.ap_ready = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_ready;
    assign module_intf_168.ap_done = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_done;
    assign module_intf_168.ap_continue = 1'b1;
    assign module_intf_168.finish = finish;
    csv_file_dump mstatus_csv_dumper_168;
    nodf_module_monitor module_monitor_168;
    nodf_module_intf module_intf_169(clock,reset);
    assign module_intf_169.ap_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_start;
    assign module_intf_169.ap_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_ready;
    assign module_intf_169.ap_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_done;
    assign module_intf_169.ap_continue = 1'b1;
    assign module_intf_169.finish = finish;
    csv_file_dump mstatus_csv_dumper_169;
    nodf_module_monitor module_monitor_169;
    nodf_module_intf module_intf_170(clock,reset);
    assign module_intf_170.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_start;
    assign module_intf_170.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ready;
    assign module_intf_170.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_done;
    assign module_intf_170.ap_continue = 1'b1;
    assign module_intf_170.finish = finish;
    csv_file_dump mstatus_csv_dumper_170;
    nodf_module_monitor module_monitor_170;
    nodf_module_intf module_intf_171(clock,reset);
    assign module_intf_171.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_start;
    assign module_intf_171.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_ready;
    assign module_intf_171.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_done;
    assign module_intf_171.ap_continue = 1'b1;
    assign module_intf_171.finish = finish;
    csv_file_dump mstatus_csv_dumper_171;
    nodf_module_monitor module_monitor_171;
    nodf_module_intf module_intf_172(clock,reset);
    assign module_intf_172.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_91_1_fu_244.ap_start;
    assign module_intf_172.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_91_1_fu_244.ap_ready;
    assign module_intf_172.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_91_1_fu_244.ap_done;
    assign module_intf_172.ap_continue = 1'b1;
    assign module_intf_172.finish = finish;
    csv_file_dump mstatus_csv_dumper_172;
    nodf_module_monitor module_monitor_172;
    nodf_module_intf module_intf_173(clock,reset);
    assign module_intf_173.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_start;
    assign module_intf_173.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_ready;
    assign module_intf_173.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_done;
    assign module_intf_173.ap_continue = 1'b1;
    assign module_intf_173.finish = finish;
    csv_file_dump mstatus_csv_dumper_173;
    nodf_module_monitor module_monitor_173;
    nodf_module_intf module_intf_174(clock,reset);
    assign module_intf_174.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_693_10_fu_260.ap_start;
    assign module_intf_174.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_693_10_fu_260.ap_ready;
    assign module_intf_174.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_693_10_fu_260.ap_done;
    assign module_intf_174.ap_continue = 1'b1;
    assign module_intf_174.finish = finish;
    csv_file_dump mstatus_csv_dumper_174;
    nodf_module_monitor module_monitor_174;
    nodf_module_intf module_intf_175(clock,reset);
    assign module_intf_175.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_start;
    assign module_intf_175.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_ready;
    assign module_intf_175.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_done;
    assign module_intf_175.ap_continue = 1'b1;
    assign module_intf_175.finish = finish;
    csv_file_dump mstatus_csv_dumper_175;
    nodf_module_monitor module_monitor_175;
    nodf_module_intf module_intf_176(clock,reset);
    assign module_intf_176.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_723_14_fu_277.ap_start;
    assign module_intf_176.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_723_14_fu_277.ap_ready;
    assign module_intf_176.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_723_14_fu_277.ap_done;
    assign module_intf_176.ap_continue = 1'b1;
    assign module_intf_176.finish = finish;
    csv_file_dump mstatus_csv_dumper_176;
    nodf_module_monitor module_monitor_176;
    nodf_module_intf module_intf_177(clock,reset);
    assign module_intf_177.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_start;
    assign module_intf_177.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_ready;
    assign module_intf_177.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_done;
    assign module_intf_177.ap_continue = 1'b1;
    assign module_intf_177.finish = finish;
    csv_file_dump mstatus_csv_dumper_177;
    nodf_module_monitor module_monitor_177;
    nodf_module_intf module_intf_178(clock,reset);
    assign module_intf_178.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_91_14_fu_296.ap_start;
    assign module_intf_178.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_91_14_fu_296.ap_ready;
    assign module_intf_178.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_91_14_fu_296.ap_done;
    assign module_intf_178.ap_continue = 1'b1;
    assign module_intf_178.finish = finish;
    csv_file_dump mstatus_csv_dumper_178;
    nodf_module_monitor module_monitor_178;
    nodf_module_intf module_intf_179(clock,reset);
    assign module_intf_179.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_start;
    assign module_intf_179.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_ready;
    assign module_intf_179.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_done;
    assign module_intf_179.ap_continue = 1'b1;
    assign module_intf_179.finish = finish;
    csv_file_dump mstatus_csv_dumper_179;
    nodf_module_monitor module_monitor_179;
    nodf_module_intf module_intf_180(clock,reset);
    assign module_intf_180.ap_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_630_6_fu_312.ap_start;
    assign module_intf_180.ap_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_630_6_fu_312.ap_ready;
    assign module_intf_180.ap_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_630_6_fu_312.ap_done;
    assign module_intf_180.ap_continue = 1'b1;
    assign module_intf_180.finish = finish;
    csv_file_dump mstatus_csv_dumper_180;
    nodf_module_monitor module_monitor_180;

    pp_loop_intf #(7) pp_loop_intf_1(clock,reset);
    assign pp_loop_intf_1.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_ST_fsm_state2;
    assign pp_loop_intf_1.pre_states_valid = 1'b1;
    assign pp_loop_intf_1.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_ST_fsm_state8;
    assign pp_loop_intf_1.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_1.post_loop_state1 = 7'h0;
    assign pp_loop_intf_1.post_states_valid[1] = 1'b0;
    assign pp_loop_intf_1.iter_start_state = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_1.iter_start_block = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.iter_end_state = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_enable_reg_pp0_iter1;
    assign pp_loop_intf_1.iter_end_block = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_1.loop_quit_state = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_1.quit_at_end = 1'b0;
    assign pp_loop_intf_1.cur_state = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.ap_CS_fsm;
    assign pp_loop_intf_1.finish = finish;
    csv_file_dump pp_loop_csv_dumper_1;
    pp_loop_monitor #(7) pp_loop_monitor_1;
    pp_loop_intf #(5) pp_loop_intf_2(clock,reset);
    assign pp_loop_intf_2.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_ST_fsm_state1;
    assign pp_loop_intf_2.pre_states_valid = 1'b1;
    assign pp_loop_intf_2.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_ST_fsm_state5;
    assign pp_loop_intf_2.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_2.post_loop_state1 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_ST_fsm_state6;
    assign pp_loop_intf_2.post_states_valid[1] = 1'b1;
    assign pp_loop_intf_2.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_2.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_2.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_2.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_2.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_enable_reg_pp0_iter1;
    assign pp_loop_intf_2.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_2.loop_quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_2.quit_at_end = 1'b1;
    assign pp_loop_intf_2.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_533_2_fu_180.ap_CS_fsm;
    assign pp_loop_intf_2.finish = finish;
    csv_file_dump pp_loop_csv_dumper_2;
    pp_loop_monitor #(5) pp_loop_monitor_2;
    pp_loop_intf #(7) pp_loop_intf_3(clock,reset);
    assign pp_loop_intf_3.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_ST_fsm_state2;
    assign pp_loop_intf_3.pre_states_valid = 1'b1;
    assign pp_loop_intf_3.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_ST_fsm_state8;
    assign pp_loop_intf_3.post_states_valid[0] = 1'b1;
    assign pp_loop_intf_3.post_loop_state1 = 7'h0;
    assign pp_loop_intf_3.post_states_valid[1] = 1'b0;
    assign pp_loop_intf_3.iter_start_state = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_3.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_enable_reg_pp0_iter0;
    assign pp_loop_intf_3.iter_start_block = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_3.iter_end_state = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_3.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_enable_reg_pp0_iter1;
    assign pp_loop_intf_3.iter_end_block = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_block_pp0_stage0_subdone;
    assign pp_loop_intf_3.loop_quit_state = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_ST_fsm_pp0_stage0;
    assign pp_loop_intf_3.quit_at_end = 1'b0;
    assign pp_loop_intf_3.cur_state = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.ap_CS_fsm;
    assign pp_loop_intf_3.finish = finish;
    csv_file_dump pp_loop_csv_dumper_3;
    pp_loop_monitor #(7) pp_loop_monitor_3;
    seq_loop_intf#(76) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state23;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state32;
    assign seq_loop_intf_1.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.post_loop_state1 = 76'h0;
    assign seq_loop_intf_1.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state24;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_dpu_keygen.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_dpu_keygen.ap_ST_fsm_state24;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state31;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(76) seq_loop_monitor_1;
    seq_loop_intf#(76) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state13;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state35;
    assign seq_loop_intf_2.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.post_loop_state1 = 76'h0;
    assign seq_loop_intf_2.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state14;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_dpu_keygen.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_dpu_keygen.ap_ST_fsm_state14;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state34;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(76) seq_loop_monitor_2;
    seq_loop_intf#(76) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state14;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state42;
    assign seq_loop_intf_3.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.post_loop_state1 = 76'h0;
    assign seq_loop_intf_3.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state35;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_dpu_keygen.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_dpu_keygen.ap_ST_fsm_state35;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state41;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(76) seq_loop_monitor_3;
    seq_loop_intf#(76) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state35;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state46;
    assign seq_loop_intf_4.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.post_loop_state1 = 76'h0;
    assign seq_loop_intf_4.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state42;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_dpu_keygen.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_dpu_keygen.ap_ST_fsm_state42;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_dpu_keygen.ap_ST_fsm_state45;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(76) seq_loop_monitor_4;
    seq_loop_intf#(198) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state1;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state198;
    assign seq_loop_intf_5.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.post_loop_state1 = 198'h0;
    assign seq_loop_intf_5.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state64;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state64;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state91;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(198) seq_loop_monitor_5;
    seq_loop_intf#(198) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state1;
    assign seq_loop_intf_6.pre_states_valid = 1'b1;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state198;
    assign seq_loop_intf_6.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.post_loop_state1 = 198'h0;
    assign seq_loop_intf_6.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state2;
    assign seq_loop_intf_6.quit_states_valid = 1'b1;
    assign seq_loop_intf_6.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state2;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state18;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(198) seq_loop_monitor_6;
    seq_loop_intf#(198) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state1;
    assign seq_loop_intf_7.pre_states_valid = 1'b1;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state198;
    assign seq_loop_intf_7.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.post_loop_state1 = 198'h0;
    assign seq_loop_intf_7.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state137;
    assign seq_loop_intf_7.quit_states_valid = 1'b1;
    assign seq_loop_intf_7.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state137;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.ap_ST_fsm_state152;
    assign seq_loop_intf_7.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(198) seq_loop_monitor_7;
    seq_loop_intf#(13) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state1;
    assign seq_loop_intf_8.pre_states_valid = 1'b1;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state3;
    assign seq_loop_intf_8.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.post_loop_state1 = 13'h0;
    assign seq_loop_intf_8.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state2;
    assign seq_loop_intf_8.quit_states_valid = 1'b1;
    assign seq_loop_intf_8.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state2;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state2;
    assign seq_loop_intf_8.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_8.one_state_loop = 1'b1;
    assign seq_loop_intf_8.one_state_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state2_blk;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(13) seq_loop_monitor_8;
    seq_loop_intf#(13) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state2;
    assign seq_loop_intf_9.pre_states_valid = 1'b1;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state7;
    assign seq_loop_intf_9.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.post_loop_state1 = 13'h0;
    assign seq_loop_intf_9.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state3;
    assign seq_loop_intf_9.quit_states_valid = 1'b1;
    assign seq_loop_intf_9.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state3;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.ap_ST_fsm_state6;
    assign seq_loop_intf_9.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(13) seq_loop_monitor_9;
    seq_loop_intf#(28) seq_loop_intf_10(clock,reset);
    assign seq_loop_intf_10.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state14;
    assign seq_loop_intf_10.pre_states_valid = 1'b1;
    assign seq_loop_intf_10.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state17;
    assign seq_loop_intf_10.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.post_loop_state1 = 28'h0;
    assign seq_loop_intf_10.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state15;
    assign seq_loop_intf_10.quit_states_valid = 1'b1;
    assign seq_loop_intf_10.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_CS_fsm;
    assign seq_loop_intf_10.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state15;
    assign seq_loop_intf_10.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state16;
    assign seq_loop_intf_10.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_10.one_state_loop = 1'b0;
    assign seq_loop_intf_10.one_state_block = 1'b0;
    assign seq_loop_intf_10.finish = finish;
    csv_file_dump seq_loop_csv_dumper_10;
    seq_loop_monitor #(28) seq_loop_monitor_10;
    seq_loop_intf#(28) seq_loop_intf_11(clock,reset);
    assign seq_loop_intf_11.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_ST_fsm_state14;
    assign seq_loop_intf_11.pre_states_valid = 1'b1;
    assign seq_loop_intf_11.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_ST_fsm_state17;
    assign seq_loop_intf_11.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.post_loop_state1 = 28'h0;
    assign seq_loop_intf_11.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_ST_fsm_state15;
    assign seq_loop_intf_11.quit_states_valid = 1'b1;
    assign seq_loop_intf_11.cur_state = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_CS_fsm;
    assign seq_loop_intf_11.iter_start_state = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_ST_fsm_state15;
    assign seq_loop_intf_11.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_2_fu_626.grp_KeccakF1600_StatePermute_fu_178.ap_ST_fsm_state16;
    assign seq_loop_intf_11.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_11.one_state_loop = 1'b0;
    assign seq_loop_intf_11.one_state_block = 1'b0;
    assign seq_loop_intf_11.finish = finish;
    csv_file_dump seq_loop_csv_dumper_11;
    seq_loop_monitor #(28) seq_loop_monitor_11;
    seq_loop_intf#(21) seq_loop_intf_12(clock,reset);
    assign seq_loop_intf_12.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state1;
    assign seq_loop_intf_12.pre_states_valid = 1'b1;
    assign seq_loop_intf_12.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state3;
    assign seq_loop_intf_12.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.post_loop_state1 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state6;
    assign seq_loop_intf_12.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_12.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state2;
    assign seq_loop_intf_12.quit_states_valid = 1'b1;
    assign seq_loop_intf_12.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_CS_fsm;
    assign seq_loop_intf_12.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state2;
    assign seq_loop_intf_12.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state2;
    assign seq_loop_intf_12.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_12.one_state_loop = 1'b1;
    assign seq_loop_intf_12.one_state_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state2_blk;
    assign seq_loop_intf_12.finish = finish;
    csv_file_dump seq_loop_csv_dumper_12;
    seq_loop_monitor #(21) seq_loop_monitor_12;
    seq_loop_intf#(21) seq_loop_intf_13(clock,reset);
    assign seq_loop_intf_13.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state10;
    assign seq_loop_intf_13.pre_states_valid = 1'b1;
    assign seq_loop_intf_13.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state15;
    assign seq_loop_intf_13.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.post_loop_state1 = 21'h0;
    assign seq_loop_intf_13.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state11;
    assign seq_loop_intf_13.quit_states_valid = 1'b1;
    assign seq_loop_intf_13.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_CS_fsm;
    assign seq_loop_intf_13.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state11;
    assign seq_loop_intf_13.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.ap_ST_fsm_state14;
    assign seq_loop_intf_13.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_13.one_state_loop = 1'b0;
    assign seq_loop_intf_13.one_state_block = 1'b0;
    assign seq_loop_intf_13.finish = finish;
    csv_file_dump seq_loop_csv_dumper_13;
    seq_loop_monitor #(21) seq_loop_monitor_13;
    seq_loop_intf#(28) seq_loop_intf_14(clock,reset);
    assign seq_loop_intf_14.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state14;
    assign seq_loop_intf_14.pre_states_valid = 1'b1;
    assign seq_loop_intf_14.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state17;
    assign seq_loop_intf_14.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.post_loop_state1 = 28'h0;
    assign seq_loop_intf_14.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state15;
    assign seq_loop_intf_14.quit_states_valid = 1'b1;
    assign seq_loop_intf_14.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_CS_fsm;
    assign seq_loop_intf_14.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state15;
    assign seq_loop_intf_14.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state16;
    assign seq_loop_intf_14.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_14.one_state_loop = 1'b0;
    assign seq_loop_intf_14.one_state_block = 1'b0;
    assign seq_loop_intf_14.finish = finish;
    csv_file_dump seq_loop_csv_dumper_14;
    seq_loop_monitor #(28) seq_loop_monitor_14;
    seq_loop_intf#(28) seq_loop_intf_15(clock,reset);
    assign seq_loop_intf_15.pre_loop_state0 = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_ST_fsm_state14;
    assign seq_loop_intf_15.pre_states_valid = 1'b1;
    assign seq_loop_intf_15.post_loop_state0 = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_ST_fsm_state17;
    assign seq_loop_intf_15.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.post_loop_state1 = 28'h0;
    assign seq_loop_intf_15.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.quit_loop_state0 = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_ST_fsm_state15;
    assign seq_loop_intf_15.quit_states_valid = 1'b1;
    assign seq_loop_intf_15.cur_state = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_CS_fsm;
    assign seq_loop_intf_15.iter_start_state = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_ST_fsm_state15;
    assign seq_loop_intf_15.iter_end_state0 = AESL_inst_dpu_keygen.grp_KeccakF1600_StatePermute_fu_650.ap_ST_fsm_state16;
    assign seq_loop_intf_15.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_15.one_state_loop = 1'b0;
    assign seq_loop_intf_15.one_state_block = 1'b0;
    assign seq_loop_intf_15.finish = finish;
    csv_file_dump seq_loop_csv_dumper_15;
    seq_loop_monitor #(28) seq_loop_monitor_15;
    seq_loop_intf#(6) seq_loop_intf_16(clock,reset);
    assign seq_loop_intf_16.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_ST_fsm_state1;
    assign seq_loop_intf_16.pre_states_valid = 1'b1;
    assign seq_loop_intf_16.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_ST_fsm_state5;
    assign seq_loop_intf_16.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.post_loop_state1 = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_ST_fsm_state6;
    assign seq_loop_intf_16.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_16.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_ST_fsm_state4;
    assign seq_loop_intf_16.quit_states_valid = 1'b1;
    assign seq_loop_intf_16.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_CS_fsm;
    assign seq_loop_intf_16.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_ST_fsm_state2;
    assign seq_loop_intf_16.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_503_2_fu_663.ap_ST_fsm_state4;
    assign seq_loop_intf_16.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_16.one_state_loop = 1'b0;
    assign seq_loop_intf_16.one_state_block = 1'b0;
    assign seq_loop_intf_16.finish = finish;
    csv_file_dump seq_loop_csv_dumper_16;
    seq_loop_monitor #(6) seq_loop_monitor_16;
    seq_loop_intf#(16) seq_loop_intf_17(clock,reset);
    assign seq_loop_intf_17.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state1;
    assign seq_loop_intf_17.pre_states_valid = 1'b1;
    assign seq_loop_intf_17.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state3;
    assign seq_loop_intf_17.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.post_loop_state1 = 16'h0;
    assign seq_loop_intf_17.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state2;
    assign seq_loop_intf_17.quit_states_valid = 1'b1;
    assign seq_loop_intf_17.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_CS_fsm;
    assign seq_loop_intf_17.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state2;
    assign seq_loop_intf_17.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state2;
    assign seq_loop_intf_17.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_17.one_state_loop = 1'b1;
    assign seq_loop_intf_17.one_state_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state2_blk;
    assign seq_loop_intf_17.finish = finish;
    csv_file_dump seq_loop_csv_dumper_17;
    seq_loop_monitor #(16) seq_loop_monitor_17;
    seq_loop_intf#(16) seq_loop_intf_18(clock,reset);
    assign seq_loop_intf_18.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state9;
    assign seq_loop_intf_18.pre_states_valid = 1'b1;
    assign seq_loop_intf_18.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state1;
    assign seq_loop_intf_18.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.post_loop_state1 = 16'h0;
    assign seq_loop_intf_18.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_18.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state10;
    assign seq_loop_intf_18.quit_states_valid = 1'b1;
    assign seq_loop_intf_18.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_CS_fsm;
    assign seq_loop_intf_18.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state10;
    assign seq_loop_intf_18.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.ap_ST_fsm_state16;
    assign seq_loop_intf_18.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_18.one_state_loop = 1'b0;
    assign seq_loop_intf_18.one_state_block = 1'b0;
    assign seq_loop_intf_18.finish = finish;
    csv_file_dump seq_loop_csv_dumper_18;
    seq_loop_monitor #(16) seq_loop_monitor_18;
    seq_loop_intf#(13) seq_loop_intf_19(clock,reset);
    assign seq_loop_intf_19.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state1;
    assign seq_loop_intf_19.pre_states_valid = 1'b1;
    assign seq_loop_intf_19.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state3;
    assign seq_loop_intf_19.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.post_loop_state1 = 13'h0;
    assign seq_loop_intf_19.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_19.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state2;
    assign seq_loop_intf_19.quit_states_valid = 1'b1;
    assign seq_loop_intf_19.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_CS_fsm;
    assign seq_loop_intf_19.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state2;
    assign seq_loop_intf_19.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state2;
    assign seq_loop_intf_19.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_19.one_state_loop = 1'b1;
    assign seq_loop_intf_19.one_state_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state2_blk;
    assign seq_loop_intf_19.finish = finish;
    csv_file_dump seq_loop_csv_dumper_19;
    seq_loop_monitor #(13) seq_loop_monitor_19;
    seq_loop_intf#(13) seq_loop_intf_20(clock,reset);
    assign seq_loop_intf_20.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state2;
    assign seq_loop_intf_20.pre_states_valid = 1'b1;
    assign seq_loop_intf_20.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state7;
    assign seq_loop_intf_20.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.post_loop_state1 = 13'h0;
    assign seq_loop_intf_20.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state3;
    assign seq_loop_intf_20.quit_states_valid = 1'b1;
    assign seq_loop_intf_20.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_CS_fsm;
    assign seq_loop_intf_20.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state3;
    assign seq_loop_intf_20.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.ap_ST_fsm_state6;
    assign seq_loop_intf_20.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_20.one_state_loop = 1'b0;
    assign seq_loop_intf_20.one_state_block = 1'b0;
    assign seq_loop_intf_20.finish = finish;
    csv_file_dump seq_loop_csv_dumper_20;
    seq_loop_monitor #(13) seq_loop_monitor_20;
    seq_loop_intf#(28) seq_loop_intf_21(clock,reset);
    assign seq_loop_intf_21.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state14;
    assign seq_loop_intf_21.pre_states_valid = 1'b1;
    assign seq_loop_intf_21.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state17;
    assign seq_loop_intf_21.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.post_loop_state1 = 28'h0;
    assign seq_loop_intf_21.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state15;
    assign seq_loop_intf_21.quit_states_valid = 1'b1;
    assign seq_loop_intf_21.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_CS_fsm;
    assign seq_loop_intf_21.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state15;
    assign seq_loop_intf_21.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_KeccakF1600_StatePermute_fu_164.ap_ST_fsm_state16;
    assign seq_loop_intf_21.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_21.one_state_loop = 1'b0;
    assign seq_loop_intf_21.one_state_block = 1'b0;
    assign seq_loop_intf_21.finish = finish;
    csv_file_dump seq_loop_csv_dumper_21;
    seq_loop_monitor #(28) seq_loop_monitor_21;
    seq_loop_intf#(21) seq_loop_intf_22(clock,reset);
    assign seq_loop_intf_22.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state1;
    assign seq_loop_intf_22.pre_states_valid = 1'b1;
    assign seq_loop_intf_22.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state3;
    assign seq_loop_intf_22.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.post_loop_state1 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state6;
    assign seq_loop_intf_22.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_22.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state2;
    assign seq_loop_intf_22.quit_states_valid = 1'b1;
    assign seq_loop_intf_22.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_CS_fsm;
    assign seq_loop_intf_22.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state2;
    assign seq_loop_intf_22.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state2;
    assign seq_loop_intf_22.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_22.one_state_loop = 1'b1;
    assign seq_loop_intf_22.one_state_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state2_blk;
    assign seq_loop_intf_22.finish = finish;
    csv_file_dump seq_loop_csv_dumper_22;
    seq_loop_monitor #(21) seq_loop_monitor_22;
    seq_loop_intf#(21) seq_loop_intf_23(clock,reset);
    assign seq_loop_intf_23.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state10;
    assign seq_loop_intf_23.pre_states_valid = 1'b1;
    assign seq_loop_intf_23.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state15;
    assign seq_loop_intf_23.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.post_loop_state1 = 21'h0;
    assign seq_loop_intf_23.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_23.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state11;
    assign seq_loop_intf_23.quit_states_valid = 1'b1;
    assign seq_loop_intf_23.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_CS_fsm;
    assign seq_loop_intf_23.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state11;
    assign seq_loop_intf_23.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.ap_ST_fsm_state14;
    assign seq_loop_intf_23.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_23.one_state_loop = 1'b0;
    assign seq_loop_intf_23.one_state_block = 1'b0;
    assign seq_loop_intf_23.finish = finish;
    csv_file_dump seq_loop_csv_dumper_23;
    seq_loop_monitor #(21) seq_loop_monitor_23;
    seq_loop_intf#(28) seq_loop_intf_24(clock,reset);
    assign seq_loop_intf_24.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state14;
    assign seq_loop_intf_24.pre_states_valid = 1'b1;
    assign seq_loop_intf_24.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state17;
    assign seq_loop_intf_24.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.post_loop_state1 = 28'h0;
    assign seq_loop_intf_24.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_24.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state15;
    assign seq_loop_intf_24.quit_states_valid = 1'b1;
    assign seq_loop_intf_24.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_CS_fsm;
    assign seq_loop_intf_24.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state15;
    assign seq_loop_intf_24.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_KeccakF1600_StatePermute_fu_265.ap_ST_fsm_state16;
    assign seq_loop_intf_24.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_24.one_state_loop = 1'b0;
    assign seq_loop_intf_24.one_state_block = 1'b0;
    assign seq_loop_intf_24.finish = finish;
    csv_file_dump seq_loop_csv_dumper_24;
    seq_loop_monitor #(28) seq_loop_monitor_24;
    seq_loop_intf#(28) seq_loop_intf_25(clock,reset);
    assign seq_loop_intf_25.pre_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_ST_fsm_state14;
    assign seq_loop_intf_25.pre_states_valid = 1'b1;
    assign seq_loop_intf_25.post_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_ST_fsm_state17;
    assign seq_loop_intf_25.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.post_loop_state1 = 28'h0;
    assign seq_loop_intf_25.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_25.quit_loop_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_ST_fsm_state15;
    assign seq_loop_intf_25.quit_states_valid = 1'b1;
    assign seq_loop_intf_25.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_CS_fsm;
    assign seq_loop_intf_25.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_ST_fsm_state15;
    assign seq_loop_intf_25.iter_end_state0 = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_KeccakF1600_StatePermute_fu_165.ap_ST_fsm_state16;
    assign seq_loop_intf_25.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_25.one_state_loop = 1'b0;
    assign seq_loop_intf_25.one_state_block = 1'b0;
    assign seq_loop_intf_25.finish = finish;
    csv_file_dump seq_loop_csv_dumper_25;
    seq_loop_monitor #(28) seq_loop_monitor_25;
    seq_loop_intf#(6) seq_loop_intf_26(clock,reset);
    assign seq_loop_intf_26.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_ST_fsm_state1;
    assign seq_loop_intf_26.pre_states_valid = 1'b1;
    assign seq_loop_intf_26.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_ST_fsm_state1;
    assign seq_loop_intf_26.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.post_loop_state1 = 6'h0;
    assign seq_loop_intf_26.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_26.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_ST_fsm_state2;
    assign seq_loop_intf_26.quit_states_valid = 1'b1;
    assign seq_loop_intf_26.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_CS_fsm;
    assign seq_loop_intf_26.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_ST_fsm_state2;
    assign seq_loop_intf_26.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.ap_ST_fsm_state6;
    assign seq_loop_intf_26.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_26.one_state_loop = 1'b0;
    assign seq_loop_intf_26.one_state_block = 1'b0;
    assign seq_loop_intf_26.finish = finish;
    csv_file_dump seq_loop_csv_dumper_26;
    seq_loop_monitor #(6) seq_loop_monitor_26;
    seq_loop_intf#(6) seq_loop_intf_27(clock,reset);
    assign seq_loop_intf_27.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_ST_fsm_state1;
    assign seq_loop_intf_27.pre_states_valid = 1'b1;
    assign seq_loop_intf_27.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_ST_fsm_state6;
    assign seq_loop_intf_27.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.post_loop_state1 = 6'h0;
    assign seq_loop_intf_27.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_27.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_ST_fsm_state2;
    assign seq_loop_intf_27.quit_states_valid = 1'b1;
    assign seq_loop_intf_27.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_CS_fsm;
    assign seq_loop_intf_27.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_ST_fsm_state2;
    assign seq_loop_intf_27.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.ap_ST_fsm_state5;
    assign seq_loop_intf_27.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_27.one_state_loop = 1'b0;
    assign seq_loop_intf_27.one_state_block = 1'b0;
    assign seq_loop_intf_27.finish = finish;
    csv_file_dump seq_loop_csv_dumper_27;
    seq_loop_monitor #(6) seq_loop_monitor_27;
    seq_loop_intf#(28) seq_loop_intf_28(clock,reset);
    assign seq_loop_intf_28.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_ST_fsm_state14;
    assign seq_loop_intf_28.pre_states_valid = 1'b1;
    assign seq_loop_intf_28.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_ST_fsm_state17;
    assign seq_loop_intf_28.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.post_loop_state1 = 28'h0;
    assign seq_loop_intf_28.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_28.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_ST_fsm_state15;
    assign seq_loop_intf_28.quit_states_valid = 1'b1;
    assign seq_loop_intf_28.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_CS_fsm;
    assign seq_loop_intf_28.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_ST_fsm_state15;
    assign seq_loop_intf_28.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_KeccakF1600_StatePermute_fu_67.ap_ST_fsm_state16;
    assign seq_loop_intf_28.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_28.one_state_loop = 1'b0;
    assign seq_loop_intf_28.one_state_block = 1'b0;
    assign seq_loop_intf_28.finish = finish;
    csv_file_dump seq_loop_csv_dumper_28;
    seq_loop_monitor #(28) seq_loop_monitor_28;
    seq_loop_intf#(28) seq_loop_intf_29(clock,reset);
    assign seq_loop_intf_29.pre_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_ST_fsm_state14;
    assign seq_loop_intf_29.pre_states_valid = 1'b1;
    assign seq_loop_intf_29.post_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_ST_fsm_state17;
    assign seq_loop_intf_29.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.post_loop_state1 = 28'h0;
    assign seq_loop_intf_29.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_29.quit_loop_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_ST_fsm_state15;
    assign seq_loop_intf_29.quit_states_valid = 1'b1;
    assign seq_loop_intf_29.cur_state = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_CS_fsm;
    assign seq_loop_intf_29.iter_start_state = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_ST_fsm_state15;
    assign seq_loop_intf_29.iter_end_state0 = AESL_inst_dpu_keygen.grp_shake_squeeze_fu_761.grp_KeccakF1600_StatePermute_fu_170.ap_ST_fsm_state16;
    assign seq_loop_intf_29.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_29.one_state_loop = 1'b0;
    assign seq_loop_intf_29.one_state_block = 1'b0;
    assign seq_loop_intf_29.finish = finish;
    csv_file_dump seq_loop_csv_dumper_29;
    seq_loop_monitor #(28) seq_loop_monitor_29;
    seq_loop_intf#(25) seq_loop_intf_30(clock,reset);
    assign seq_loop_intf_30.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state1;
    assign seq_loop_intf_30.pre_states_valid = 1'b1;
    assign seq_loop_intf_30.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state25;
    assign seq_loop_intf_30.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.post_loop_state1 = 25'h0;
    assign seq_loop_intf_30.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_30.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state20;
    assign seq_loop_intf_30.quit_states_valid = 1'b1;
    assign seq_loop_intf_30.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_CS_fsm;
    assign seq_loop_intf_30.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state20;
    assign seq_loop_intf_30.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state24;
    assign seq_loop_intf_30.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_30.one_state_loop = 1'b0;
    assign seq_loop_intf_30.one_state_block = 1'b0;
    assign seq_loop_intf_30.finish = finish;
    csv_file_dump seq_loop_csv_dumper_30;
    seq_loop_monitor #(25) seq_loop_monitor_30;
    seq_loop_intf#(25) seq_loop_intf_31(clock,reset);
    assign seq_loop_intf_31.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state1;
    assign seq_loop_intf_31.pre_states_valid = 1'b1;
    assign seq_loop_intf_31.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state25;
    assign seq_loop_intf_31.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.post_loop_state1 = 25'h0;
    assign seq_loop_intf_31.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_31.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state2;
    assign seq_loop_intf_31.quit_states_valid = 1'b1;
    assign seq_loop_intf_31.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_CS_fsm;
    assign seq_loop_intf_31.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state2;
    assign seq_loop_intf_31.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state5;
    assign seq_loop_intf_31.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_31.one_state_loop = 1'b0;
    assign seq_loop_intf_31.one_state_block = 1'b0;
    assign seq_loop_intf_31.finish = finish;
    csv_file_dump seq_loop_csv_dumper_31;
    seq_loop_monitor #(25) seq_loop_monitor_31;
    seq_loop_intf#(25) seq_loop_intf_32(clock,reset);
    assign seq_loop_intf_32.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state1;
    assign seq_loop_intf_32.pre_states_valid = 1'b1;
    assign seq_loop_intf_32.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state25;
    assign seq_loop_intf_32.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.post_loop_state1 = 25'h0;
    assign seq_loop_intf_32.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_32.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state6;
    assign seq_loop_intf_32.quit_states_valid = 1'b1;
    assign seq_loop_intf_32.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_CS_fsm;
    assign seq_loop_intf_32.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state6;
    assign seq_loop_intf_32.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state10;
    assign seq_loop_intf_32.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_32.one_state_loop = 1'b0;
    assign seq_loop_intf_32.one_state_block = 1'b0;
    assign seq_loop_intf_32.finish = finish;
    csv_file_dump seq_loop_csv_dumper_32;
    seq_loop_monitor #(25) seq_loop_monitor_32;
    seq_loop_intf#(25) seq_loop_intf_33(clock,reset);
    assign seq_loop_intf_33.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state1;
    assign seq_loop_intf_33.pre_states_valid = 1'b1;
    assign seq_loop_intf_33.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state25;
    assign seq_loop_intf_33.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.post_loop_state1 = 25'h0;
    assign seq_loop_intf_33.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_33.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state16;
    assign seq_loop_intf_33.quit_states_valid = 1'b1;
    assign seq_loop_intf_33.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_CS_fsm;
    assign seq_loop_intf_33.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state16;
    assign seq_loop_intf_33.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state19;
    assign seq_loop_intf_33.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_33.one_state_loop = 1'b0;
    assign seq_loop_intf_33.one_state_block = 1'b0;
    assign seq_loop_intf_33.finish = finish;
    csv_file_dump seq_loop_csv_dumper_33;
    seq_loop_monitor #(25) seq_loop_monitor_33;
    seq_loop_intf#(25) seq_loop_intf_34(clock,reset);
    assign seq_loop_intf_34.pre_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state1;
    assign seq_loop_intf_34.pre_states_valid = 1'b1;
    assign seq_loop_intf_34.post_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state25;
    assign seq_loop_intf_34.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.post_loop_state1 = 25'h0;
    assign seq_loop_intf_34.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_34.quit_loop_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state11;
    assign seq_loop_intf_34.quit_states_valid = 1'b1;
    assign seq_loop_intf_34.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_CS_fsm;
    assign seq_loop_intf_34.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state11;
    assign seq_loop_intf_34.iter_end_state0 = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.ap_ST_fsm_state15;
    assign seq_loop_intf_34.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_34.one_state_loop = 1'b0;
    assign seq_loop_intf_34.one_state_block = 1'b0;
    assign seq_loop_intf_34.finish = finish;
    csv_file_dump seq_loop_csv_dumper_34;
    seq_loop_monitor #(25) seq_loop_monitor_34;
    upc_loop_intf#(32) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_1.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_POW2ROUND_LOOP1_fu_715.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b0;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(32) upc_loop_monitor_1;
    upc_loop_intf#(31) upc_loop_intf_2(clock,reset);
    assign upc_loop_intf_2.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_CS_fsm;
    assign upc_loop_intf_2.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_2.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_2.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_2.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_2.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_start;
    assign upc_loop_intf_2.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_ready;
    assign upc_loop_intf_2.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_CADDQ_LOOP1_fu_737.ap_done_int;
    assign upc_loop_intf_2.loop_continue = 1'b1;
    assign upc_loop_intf_2.quit_at_end = 1'b0;
    assign upc_loop_intf_2.finish = finish;
    csv_file_dump upc_loop_csv_dumper_2;
    upc_loop_monitor #(31) upc_loop_monitor_2;
    upc_loop_intf#(34) upc_loop_intf_3(clock,reset);
    assign upc_loop_intf_3.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_CS_fsm;
    assign upc_loop_intf_3.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_3.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_3.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_3.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_3.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_start;
    assign upc_loop_intf_3.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_ready;
    assign upc_loop_intf_3.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP1_fu_757.ap_done_int;
    assign upc_loop_intf_3.loop_continue = 1'b1;
    assign upc_loop_intf_3.quit_at_end = 1'b0;
    assign upc_loop_intf_3.finish = finish;
    csv_file_dump upc_loop_csv_dumper_3;
    upc_loop_monitor #(34) upc_loop_monitor_3;
    upc_loop_intf#(31) upc_loop_intf_4(clock,reset);
    assign upc_loop_intf_4.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_CS_fsm;
    assign upc_loop_intf_4.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_4.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_4.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_4.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_4.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_start;
    assign upc_loop_intf_4.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_ready;
    assign upc_loop_intf_4.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP1_fu_776.ap_done_int;
    assign upc_loop_intf_4.loop_continue = 1'b1;
    assign upc_loop_intf_4.quit_at_end = 1'b0;
    assign upc_loop_intf_4.finish = finish;
    csv_file_dump upc_loop_csv_dumper_4;
    upc_loop_monitor #(31) upc_loop_monitor_4;
    upc_loop_intf#(33) upc_loop_intf_5(clock,reset);
    assign upc_loop_intf_5.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_CS_fsm;
    assign upc_loop_intf_5.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_5.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_5.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_5.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_5.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_start;
    assign upc_loop_intf_5.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_ready;
    assign upc_loop_intf_5.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_SUB_LOOP1_fu_796.ap_done_int;
    assign upc_loop_intf_5.loop_continue = 1'b1;
    assign upc_loop_intf_5.quit_at_end = 1'b0;
    assign upc_loop_intf_5.finish = finish;
    csv_file_dump upc_loop_csv_dumper_5;
    upc_loop_monitor #(33) upc_loop_monitor_5;
    upc_loop_intf#(33) upc_loop_intf_6(clock,reset);
    assign upc_loop_intf_6.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_CS_fsm;
    assign upc_loop_intf_6.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_6.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_6.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_6.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_6.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_start;
    assign upc_loop_intf_6.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_ready;
    assign upc_loop_intf_6.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_ADD_LOOP1_fu_819.ap_done_int;
    assign upc_loop_intf_6.loop_continue = 1'b1;
    assign upc_loop_intf_6.quit_at_end = 1'b0;
    assign upc_loop_intf_6.finish = finish;
    csv_file_dump upc_loop_csv_dumper_6;
    upc_loop_monitor #(33) upc_loop_monitor_6;
    upc_loop_intf#(32) upc_loop_intf_7(clock,reset);
    assign upc_loop_intf_7.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_CS_fsm;
    assign upc_loop_intf_7.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_7.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_7.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_7.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_7.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_start;
    assign upc_loop_intf_7.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_ready;
    assign upc_loop_intf_7.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP1_fu_842.ap_done_int;
    assign upc_loop_intf_7.loop_continue = 1'b1;
    assign upc_loop_intf_7.quit_at_end = 1'b0;
    assign upc_loop_intf_7.finish = finish;
    csv_file_dump upc_loop_csv_dumper_7;
    upc_loop_monitor #(32) upc_loop_monitor_7;
    upc_loop_intf#(31) upc_loop_intf_8(clock,reset);
    assign upc_loop_intf_8.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_CS_fsm;
    assign upc_loop_intf_8.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_8.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_8.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_8.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_8.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_start;
    assign upc_loop_intf_8.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_ready;
    assign upc_loop_intf_8.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP2_fu_857.ap_done_int;
    assign upc_loop_intf_8.loop_continue = 1'b1;
    assign upc_loop_intf_8.quit_at_end = 1'b0;
    assign upc_loop_intf_8.finish = finish;
    csv_file_dump upc_loop_csv_dumper_8;
    upc_loop_monitor #(31) upc_loop_monitor_8;
    upc_loop_intf#(31) upc_loop_intf_9(clock,reset);
    assign upc_loop_intf_9.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_CS_fsm;
    assign upc_loop_intf_9.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_9.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_9.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_9.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_9.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_start;
    assign upc_loop_intf_9.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_ready;
    assign upc_loop_intf_9.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP3_fu_871.ap_done_int;
    assign upc_loop_intf_9.loop_continue = 1'b1;
    assign upc_loop_intf_9.quit_at_end = 1'b0;
    assign upc_loop_intf_9.finish = finish;
    csv_file_dump upc_loop_csv_dumper_9;
    upc_loop_monitor #(31) upc_loop_monitor_9;
    upc_loop_intf#(33) upc_loop_intf_10(clock,reset);
    assign upc_loop_intf_10.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_CS_fsm;
    assign upc_loop_intf_10.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_10.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_10.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_10.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_10.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_start;
    assign upc_loop_intf_10.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_ready;
    assign upc_loop_intf_10.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP4_fu_885.ap_done_int;
    assign upc_loop_intf_10.loop_continue = 1'b1;
    assign upc_loop_intf_10.quit_at_end = 1'b0;
    assign upc_loop_intf_10.finish = finish;
    csv_file_dump upc_loop_csv_dumper_10;
    upc_loop_monitor #(33) upc_loop_monitor_10;
    upc_loop_intf#(31) upc_loop_intf_11(clock,reset);
    assign upc_loop_intf_11.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_CS_fsm;
    assign upc_loop_intf_11.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_11.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_11.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_11.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_11.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_start;
    assign upc_loop_intf_11.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_ready;
    assign upc_loop_intf_11.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_NTT_LOOP5_fu_901.ap_done_int;
    assign upc_loop_intf_11.loop_continue = 1'b1;
    assign upc_loop_intf_11.quit_at_end = 1'b0;
    assign upc_loop_intf_11.finish = finish;
    csv_file_dump upc_loop_csv_dumper_11;
    upc_loop_monitor #(31) upc_loop_monitor_11;
    upc_loop_intf#(34) upc_loop_intf_12(clock,reset);
    assign upc_loop_intf_12.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_CS_fsm;
    assign upc_loop_intf_12.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_12.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_12.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_12.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_12.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_start;
    assign upc_loop_intf_12.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_ready;
    assign upc_loop_intf_12.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP1_fu_917.ap_done_int;
    assign upc_loop_intf_12.loop_continue = 1'b1;
    assign upc_loop_intf_12.quit_at_end = 1'b0;
    assign upc_loop_intf_12.finish = finish;
    csv_file_dump upc_loop_csv_dumper_12;
    upc_loop_monitor #(34) upc_loop_monitor_12;
    upc_loop_intf#(31) upc_loop_intf_13(clock,reset);
    assign upc_loop_intf_13.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_CS_fsm;
    assign upc_loop_intf_13.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_13.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_13.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_13.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_13.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_start;
    assign upc_loop_intf_13.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_ready;
    assign upc_loop_intf_13.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP2_fu_933.ap_done_int;
    assign upc_loop_intf_13.loop_continue = 1'b1;
    assign upc_loop_intf_13.quit_at_end = 1'b0;
    assign upc_loop_intf_13.finish = finish;
    csv_file_dump upc_loop_csv_dumper_13;
    upc_loop_monitor #(31) upc_loop_monitor_13;
    upc_loop_intf#(31) upc_loop_intf_14(clock,reset);
    assign upc_loop_intf_14.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_CS_fsm;
    assign upc_loop_intf_14.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_14.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_14.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_14.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_14.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_14.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_start;
    assign upc_loop_intf_14.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_ready;
    assign upc_loop_intf_14.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP3_fu_947.ap_done_int;
    assign upc_loop_intf_14.loop_continue = 1'b1;
    assign upc_loop_intf_14.quit_at_end = 1'b0;
    assign upc_loop_intf_14.finish = finish;
    csv_file_dump upc_loop_csv_dumper_14;
    upc_loop_monitor #(31) upc_loop_monitor_14;
    upc_loop_intf#(33) upc_loop_intf_15(clock,reset);
    assign upc_loop_intf_15.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_CS_fsm;
    assign upc_loop_intf_15.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_15.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_15.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_15.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_15.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_start;
    assign upc_loop_intf_15.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_ready;
    assign upc_loop_intf_15.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP4_fu_961.ap_done_int;
    assign upc_loop_intf_15.loop_continue = 1'b1;
    assign upc_loop_intf_15.quit_at_end = 1'b0;
    assign upc_loop_intf_15.finish = finish;
    csv_file_dump upc_loop_csv_dumper_15;
    upc_loop_monitor #(33) upc_loop_monitor_15;
    upc_loop_intf#(34) upc_loop_intf_16(clock,reset);
    assign upc_loop_intf_16.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_CS_fsm;
    assign upc_loop_intf_16.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_16.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_16.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_16.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_16.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_16.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_16.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_start;
    assign upc_loop_intf_16.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_ready;
    assign upc_loop_intf_16.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MATMUL_LOOP5_fu_976.ap_done_int;
    assign upc_loop_intf_16.loop_continue = 1'b1;
    assign upc_loop_intf_16.quit_at_end = 1'b0;
    assign upc_loop_intf_16.finish = finish;
    csv_file_dump upc_loop_csv_dumper_16;
    upc_loop_monitor #(34) upc_loop_monitor_16;
    upc_loop_intf#(31) upc_loop_intf_17(clock,reset);
    assign upc_loop_intf_17.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_CS_fsm;
    assign upc_loop_intf_17.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_17.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_17.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_17.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_17.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_start;
    assign upc_loop_intf_17.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_ready;
    assign upc_loop_intf_17.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP2_fu_992.ap_done_int;
    assign upc_loop_intf_17.loop_continue = 1'b1;
    assign upc_loop_intf_17.quit_at_end = 1'b0;
    assign upc_loop_intf_17.finish = finish;
    csv_file_dump upc_loop_csv_dumper_17;
    upc_loop_monitor #(31) upc_loop_monitor_17;
    upc_loop_intf#(31) upc_loop_intf_18(clock,reset);
    assign upc_loop_intf_18.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_CS_fsm;
    assign upc_loop_intf_18.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_18.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_18.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_18.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_18.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_start;
    assign upc_loop_intf_18.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_ready;
    assign upc_loop_intf_18.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP3_fu_1006.ap_done_int;
    assign upc_loop_intf_18.loop_continue = 1'b1;
    assign upc_loop_intf_18.quit_at_end = 1'b0;
    assign upc_loop_intf_18.finish = finish;
    csv_file_dump upc_loop_csv_dumper_18;
    upc_loop_monitor #(31) upc_loop_monitor_18;
    upc_loop_intf#(33) upc_loop_intf_19(clock,reset);
    assign upc_loop_intf_19.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_CS_fsm;
    assign upc_loop_intf_19.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_19.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_19.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_19.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_19.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_start;
    assign upc_loop_intf_19.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_ready;
    assign upc_loop_intf_19.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_MONTMUL_LOOP4_fu_1020.ap_done_int;
    assign upc_loop_intf_19.loop_continue = 1'b1;
    assign upc_loop_intf_19.quit_at_end = 1'b0;
    assign upc_loop_intf_19.finish = finish;
    csv_file_dump upc_loop_csv_dumper_19;
    upc_loop_monitor #(33) upc_loop_monitor_19;
    upc_loop_intf#(31) upc_loop_intf_20(clock,reset);
    assign upc_loop_intf_20.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_CS_fsm;
    assign upc_loop_intf_20.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_20.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_20.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_20.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_20.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_20.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_start;
    assign upc_loop_intf_20.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_ready;
    assign upc_loop_intf_20.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP2_fu_1036.ap_done_int;
    assign upc_loop_intf_20.loop_continue = 1'b1;
    assign upc_loop_intf_20.quit_at_end = 1'b0;
    assign upc_loop_intf_20.finish = finish;
    csv_file_dump upc_loop_csv_dumper_20;
    upc_loop_monitor #(31) upc_loop_monitor_20;
    upc_loop_intf#(33) upc_loop_intf_21(clock,reset);
    assign upc_loop_intf_21.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_CS_fsm;
    assign upc_loop_intf_21.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_21.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_21.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_21.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_21.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_start;
    assign upc_loop_intf_21.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_ready;
    assign upc_loop_intf_21.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_RD_LOOP3_fu_1050.ap_done_int;
    assign upc_loop_intf_21.loop_continue = 1'b1;
    assign upc_loop_intf_21.quit_at_end = 1'b0;
    assign upc_loop_intf_21.finish = finish;
    csv_file_dump upc_loop_csv_dumper_21;
    upc_loop_monitor #(33) upc_loop_monitor_21;
    upc_loop_intf#(31) upc_loop_intf_22(clock,reset);
    assign upc_loop_intf_22.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_CS_fsm;
    assign upc_loop_intf_22.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_22.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_22.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_22.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_22.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_22.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_start;
    assign upc_loop_intf_22.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_ready;
    assign upc_loop_intf_22.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP1_fu_1066.ap_done_int;
    assign upc_loop_intf_22.loop_continue = 1'b1;
    assign upc_loop_intf_22.quit_at_end = 1'b0;
    assign upc_loop_intf_22.finish = finish;
    csv_file_dump upc_loop_csv_dumper_22;
    upc_loop_monitor #(31) upc_loop_monitor_22;
    upc_loop_intf#(32) upc_loop_intf_23(clock,reset);
    assign upc_loop_intf_23.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_CS_fsm;
    assign upc_loop_intf_23.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_23.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_23.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_23.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_23.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_23.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_start;
    assign upc_loop_intf_23.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_ready;
    assign upc_loop_intf_23.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP2_fu_1080.ap_done_int;
    assign upc_loop_intf_23.loop_continue = 1'b1;
    assign upc_loop_intf_23.quit_at_end = 1'b0;
    assign upc_loop_intf_23.finish = finish;
    csv_file_dump upc_loop_csv_dumper_23;
    upc_loop_monitor #(32) upc_loop_monitor_23;
    upc_loop_intf#(31) upc_loop_intf_24(clock,reset);
    assign upc_loop_intf_24.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_CS_fsm;
    assign upc_loop_intf_24.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_24.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_24.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_24.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_24.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_24.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_start;
    assign upc_loop_intf_24.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_ready;
    assign upc_loop_intf_24.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP3_fu_1095.ap_done_int;
    assign upc_loop_intf_24.loop_continue = 1'b1;
    assign upc_loop_intf_24.quit_at_end = 1'b0;
    assign upc_loop_intf_24.finish = finish;
    csv_file_dump upc_loop_csv_dumper_24;
    upc_loop_monitor #(31) upc_loop_monitor_24;
    upc_loop_intf#(31) upc_loop_intf_25(clock,reset);
    assign upc_loop_intf_25.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_CS_fsm;
    assign upc_loop_intf_25.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_25.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_25.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_25.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_25.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_25.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_start;
    assign upc_loop_intf_25.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_ready;
    assign upc_loop_intf_25.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP4_fu_1109.ap_done_int;
    assign upc_loop_intf_25.loop_continue = 1'b1;
    assign upc_loop_intf_25.quit_at_end = 1'b0;
    assign upc_loop_intf_25.finish = finish;
    csv_file_dump upc_loop_csv_dumper_25;
    upc_loop_monitor #(31) upc_loop_monitor_25;
    upc_loop_intf#(33) upc_loop_intf_26(clock,reset);
    assign upc_loop_intf_26.cur_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_CS_fsm;
    assign upc_loop_intf_26.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.quit_state = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_26.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.quit_block = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_26.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_26.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_26.quit_enable = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_26.loop_start = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_start;
    assign upc_loop_intf_26.loop_ready = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_ready;
    assign upc_loop_intf_26.loop_done = AESL_inst_dpu_keygen.grp_dpu_func_fu_460.grp_dpu_func_Pipeline_FUNC_INTT_LOOP5_fu_1123.ap_done_int;
    assign upc_loop_intf_26.loop_continue = 1'b1;
    assign upc_loop_intf_26.quit_at_end = 1'b0;
    assign upc_loop_intf_26.finish = finish;
    csv_file_dump upc_loop_csv_dumper_26;
    upc_loop_monitor #(33) upc_loop_monitor_26;
    upc_loop_intf#(1) upc_loop_intf_27(clock,reset);
    assign upc_loop_intf_27.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_CS_fsm;
    assign upc_loop_intf_27.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_27.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_27.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_27.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_27.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_27.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_start;
    assign upc_loop_intf_27.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_ready;
    assign upc_loop_intf_27.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_42_3_VITIS_LOOP_43_4_fu_578.ap_done_int;
    assign upc_loop_intf_27.loop_continue = 1'b1;
    assign upc_loop_intf_27.quit_at_end = 1'b0;
    assign upc_loop_intf_27.finish = finish;
    csv_file_dump upc_loop_csv_dumper_27;
    upc_loop_monitor #(1) upc_loop_monitor_27;
    upc_loop_intf#(4) upc_loop_intf_28(clock,reset);
    assign upc_loop_intf_28.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_CS_fsm;
    assign upc_loop_intf_28.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_28.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_28.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_28.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_28.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_28.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_start;
    assign upc_loop_intf_28.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ready;
    assign upc_loop_intf_28.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_done_int;
    assign upc_loop_intf_28.loop_continue = 1'b1;
    assign upc_loop_intf_28.quit_at_end = 1'b0;
    assign upc_loop_intf_28.finish = finish;
    csv_file_dump upc_loop_csv_dumper_28;
    upc_loop_monitor #(4) upc_loop_monitor_28;
    upc_loop_intf#(4) upc_loop_intf_29(clock,reset);
    assign upc_loop_intf_29.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_CS_fsm;
    assign upc_loop_intf_29.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_29.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_29.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_29.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_29.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_29.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_start;
    assign upc_loop_intf_29.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ready;
    assign upc_loop_intf_29.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_done_int;
    assign upc_loop_intf_29.loop_continue = 1'b1;
    assign upc_loop_intf_29.quit_at_end = 1'b0;
    assign upc_loop_intf_29.finish = finish;
    csv_file_dump upc_loop_csv_dumper_29;
    upc_loop_monitor #(4) upc_loop_monitor_29;
    upc_loop_intf#(1) upc_loop_intf_30(clock,reset);
    assign upc_loop_intf_30.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_CS_fsm;
    assign upc_loop_intf_30.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_30.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_30.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_30.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_30.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_30.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_start;
    assign upc_loop_intf_30.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ready;
    assign upc_loop_intf_30.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_done_int;
    assign upc_loop_intf_30.loop_continue = 1'b1;
    assign upc_loop_intf_30.quit_at_end = 1'b0;
    assign upc_loop_intf_30.finish = finish;
    csv_file_dump upc_loop_csv_dumper_30;
    upc_loop_monitor #(1) upc_loop_monitor_30;
    upc_loop_intf#(1) upc_loop_intf_31(clock,reset);
    assign upc_loop_intf_31.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_CS_fsm;
    assign upc_loop_intf_31.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_31.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_31.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_31.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_31.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_31.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_start;
    assign upc_loop_intf_31.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ready;
    assign upc_loop_intf_31.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_1_fu_585.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_done_int;
    assign upc_loop_intf_31.loop_continue = 1'b1;
    assign upc_loop_intf_31.quit_at_end = 1'b0;
    assign upc_loop_intf_31.finish = finish;
    csv_file_dump upc_loop_csv_dumper_31;
    upc_loop_monitor #(1) upc_loop_monitor_31;
    upc_loop_intf#(1) upc_loop_intf_32(clock,reset);
    assign upc_loop_intf_32.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_CS_fsm;
    assign upc_loop_intf_32.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_32.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_32.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_32.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_32.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_32.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_32.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_32.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_32.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_32.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_start;
    assign upc_loop_intf_32.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_ready;
    assign upc_loop_intf_32.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_48_5_VITIS_LOOP_49_6_fu_599.ap_done_int;
    assign upc_loop_intf_32.loop_continue = 1'b1;
    assign upc_loop_intf_32.quit_at_end = 1'b0;
    assign upc_loop_intf_32.finish = finish;
    csv_file_dump upc_loop_csv_dumper_32;
    upc_loop_monitor #(1) upc_loop_monitor_32;
    upc_loop_intf#(1) upc_loop_intf_33(clock,reset);
    assign upc_loop_intf_33.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_CS_fsm;
    assign upc_loop_intf_33.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_33.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_33.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_33.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_33.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_33.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_start;
    assign upc_loop_intf_33.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_ready;
    assign upc_loop_intf_33.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_54_7_fu_606.ap_done_int;
    assign upc_loop_intf_33.loop_continue = 1'b1;
    assign upc_loop_intf_33.quit_at_end = 1'b1;
    assign upc_loop_intf_33.finish = finish;
    csv_file_dump upc_loop_csv_dumper_33;
    upc_loop_monitor #(1) upc_loop_monitor_33;
    upc_loop_intf#(1) upc_loop_intf_34(clock,reset);
    assign upc_loop_intf_34.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_CS_fsm;
    assign upc_loop_intf_34.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_34.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_34.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_34.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_34.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_34.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_34.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_34.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_34.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_34.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_start;
    assign upc_loop_intf_34.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_ready;
    assign upc_loop_intf_34.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_8_fu_612.ap_done_int;
    assign upc_loop_intf_34.loop_continue = 1'b1;
    assign upc_loop_intf_34.quit_at_end = 1'b1;
    assign upc_loop_intf_34.finish = finish;
    csv_file_dump upc_loop_csv_dumper_34;
    upc_loop_monitor #(1) upc_loop_monitor_34;
    upc_loop_intf#(1) upc_loop_intf_35(clock,reset);
    assign upc_loop_intf_35.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_CS_fsm;
    assign upc_loop_intf_35.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_35.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_35.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_35.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_35.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_35.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_35.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_35.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_35.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_35.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_start;
    assign upc_loop_intf_35.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_ready;
    assign upc_loop_intf_35.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_56_9_fu_619.ap_done_int;
    assign upc_loop_intf_35.loop_continue = 1'b1;
    assign upc_loop_intf_35.quit_at_end = 1'b1;
    assign upc_loop_intf_35.finish = finish;
    csv_file_dump upc_loop_csv_dumper_35;
    upc_loop_monitor #(1) upc_loop_monitor_35;
    upc_loop_intf#(1) upc_loop_intf_36(clock,reset);
    assign upc_loop_intf_36.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_CS_fsm;
    assign upc_loop_intf_36.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_36.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_36.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_36.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_36.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_36.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_36.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_36.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_36.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_36.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_start;
    assign upc_loop_intf_36.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ready;
    assign upc_loop_intf_36.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_done_int;
    assign upc_loop_intf_36.loop_continue = 1'b1;
    assign upc_loop_intf_36.quit_at_end = 1'b1;
    assign upc_loop_intf_36.finish = finish;
    csv_file_dump upc_loop_csv_dumper_36;
    upc_loop_monitor #(1) upc_loop_monitor_36;
    upc_loop_intf#(1) upc_loop_intf_37(clock,reset);
    assign upc_loop_intf_37.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_CS_fsm;
    assign upc_loop_intf_37.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_37.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_37.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_37.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_37.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_37.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_37.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_37.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_37.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_37.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_start;
    assign upc_loop_intf_37.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ready;
    assign upc_loop_intf_37.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_done_int;
    assign upc_loop_intf_37.loop_continue = 1'b1;
    assign upc_loop_intf_37.quit_at_end = 1'b0;
    assign upc_loop_intf_37.finish = finish;
    csv_file_dump upc_loop_csv_dumper_37;
    upc_loop_monitor #(1) upc_loop_monitor_37;
    upc_loop_intf#(1) upc_loop_intf_38(clock,reset);
    assign upc_loop_intf_38.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_CS_fsm;
    assign upc_loop_intf_38.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_38.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_38.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_38.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_38.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_38.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_38.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_38.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_38.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_38.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_start;
    assign upc_loop_intf_38.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ready;
    assign upc_loop_intf_38.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_done_int;
    assign upc_loop_intf_38.loop_continue = 1'b1;
    assign upc_loop_intf_38.quit_at_end = 1'b0;
    assign upc_loop_intf_38.finish = finish;
    csv_file_dump upc_loop_csv_dumper_38;
    upc_loop_monitor #(1) upc_loop_monitor_38;
    upc_loop_intf#(1) upc_loop_intf_39(clock,reset);
    assign upc_loop_intf_39.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_CS_fsm;
    assign upc_loop_intf_39.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_39.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_39.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_39.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_39.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_39.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_39.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_39.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_39.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_39.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_start;
    assign upc_loop_intf_39.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ready;
    assign upc_loop_intf_39.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_done_int;
    assign upc_loop_intf_39.loop_continue = 1'b1;
    assign upc_loop_intf_39.quit_at_end = 1'b0;
    assign upc_loop_intf_39.finish = finish;
    csv_file_dump upc_loop_csv_dumper_39;
    upc_loop_monitor #(1) upc_loop_monitor_39;
    upc_loop_intf#(1) upc_loop_intf_40(clock,reset);
    assign upc_loop_intf_40.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_CS_fsm;
    assign upc_loop_intf_40.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_40.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_40.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_40.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_40.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_40.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_40.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_40.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_40.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_40.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_start;
    assign upc_loop_intf_40.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ready;
    assign upc_loop_intf_40.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_done_int;
    assign upc_loop_intf_40.loop_continue = 1'b1;
    assign upc_loop_intf_40.quit_at_end = 1'b0;
    assign upc_loop_intf_40.finish = finish;
    csv_file_dump upc_loop_csv_dumper_40;
    upc_loop_monitor #(1) upc_loop_monitor_40;
    upc_loop_intf#(1) upc_loop_intf_41(clock,reset);
    assign upc_loop_intf_41.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_CS_fsm;
    assign upc_loop_intf_41.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_41.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_41.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_41.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_41.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_41.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_41.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_41.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_41.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_41.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_start;
    assign upc_loop_intf_41.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ready;
    assign upc_loop_intf_41.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_fu_640.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_done_int;
    assign upc_loop_intf_41.loop_continue = 1'b1;
    assign upc_loop_intf_41.quit_at_end = 1'b0;
    assign upc_loop_intf_41.finish = finish;
    csv_file_dump upc_loop_csv_dumper_41;
    upc_loop_monitor #(1) upc_loop_monitor_41;
    upc_loop_intf#(4) upc_loop_intf_42(clock,reset);
    assign upc_loop_intf_42.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_CS_fsm;
    assign upc_loop_intf_42.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_42.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_42.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_42.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_42.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_42.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_42.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_42.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_42.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_42.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_start;
    assign upc_loop_intf_42.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_ready;
    assign upc_loop_intf_42.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_417_2_fu_657.ap_done_int;
    assign upc_loop_intf_42.loop_continue = 1'b1;
    assign upc_loop_intf_42.quit_at_end = 1'b0;
    assign upc_loop_intf_42.finish = finish;
    csv_file_dump upc_loop_csv_dumper_42;
    upc_loop_monitor #(4) upc_loop_monitor_42;
    upc_loop_intf#(1) upc_loop_intf_43(clock,reset);
    assign upc_loop_intf_43.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_CS_fsm;
    assign upc_loop_intf_43.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_43.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_43.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_43.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_43.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_43.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_43.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_43.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_43.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_43.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_start;
    assign upc_loop_intf_43.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_ready;
    assign upc_loop_intf_43.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_1_fu_671.ap_done_int;
    assign upc_loop_intf_43.loop_continue = 1'b1;
    assign upc_loop_intf_43.quit_at_end = 1'b0;
    assign upc_loop_intf_43.finish = finish;
    csv_file_dump upc_loop_csv_dumper_43;
    upc_loop_monitor #(1) upc_loop_monitor_43;
    upc_loop_intf#(4) upc_loop_intf_44(clock,reset);
    assign upc_loop_intf_44.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_CS_fsm;
    assign upc_loop_intf_44.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_44.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_44.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_44.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_44.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_44.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_44.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_44.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_44.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_44.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_start;
    assign upc_loop_intf_44.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_ready;
    assign upc_loop_intf_44.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_369_4_fu_143.ap_done_int;
    assign upc_loop_intf_44.loop_continue = 1'b1;
    assign upc_loop_intf_44.quit_at_end = 1'b0;
    assign upc_loop_intf_44.finish = finish;
    csv_file_dump upc_loop_csv_dumper_44;
    upc_loop_monitor #(4) upc_loop_monitor_44;
    upc_loop_intf#(4) upc_loop_intf_45(clock,reset);
    assign upc_loop_intf_45.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_CS_fsm;
    assign upc_loop_intf_45.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_45.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_45.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_45.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_45.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_45.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_45.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_45.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_45.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_45.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_start;
    assign upc_loop_intf_45.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_ready;
    assign upc_loop_intf_45.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_376_5_fu_154.ap_done_int;
    assign upc_loop_intf_45.loop_continue = 1'b1;
    assign upc_loop_intf_45.quit_at_end = 1'b0;
    assign upc_loop_intf_45.finish = finish;
    csv_file_dump upc_loop_csv_dumper_45;
    upc_loop_monitor #(4) upc_loop_monitor_45;
    upc_loop_intf#(1) upc_loop_intf_46(clock,reset);
    assign upc_loop_intf_46.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_CS_fsm;
    assign upc_loop_intf_46.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_46.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_46.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_46.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_46.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_46.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_46.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_46.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_46.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_46.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_start;
    assign upc_loop_intf_46.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_ready;
    assign upc_loop_intf_46.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_385_7_fu_177.ap_done_int;
    assign upc_loop_intf_46.loop_continue = 1'b1;
    assign upc_loop_intf_46.quit_at_end = 1'b0;
    assign upc_loop_intf_46.finish = finish;
    csv_file_dump upc_loop_csv_dumper_46;
    upc_loop_monitor #(1) upc_loop_monitor_46;
    upc_loop_intf#(1) upc_loop_intf_47(clock,reset);
    assign upc_loop_intf_47.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_CS_fsm;
    assign upc_loop_intf_47.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_47.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_47.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_47.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_47.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_47.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_47.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_47.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_47.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_47.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_start;
    assign upc_loop_intf_47.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_ready;
    assign upc_loop_intf_47.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_1_fu_139.grp_shake_absorb_1_Pipeline_VITIS_LOOP_12_1_fu_187.ap_done_int;
    assign upc_loop_intf_47.loop_continue = 1'b1;
    assign upc_loop_intf_47.quit_at_end = 1'b0;
    assign upc_loop_intf_47.finish = finish;
    csv_file_dump upc_loop_csv_dumper_47;
    upc_loop_monitor #(1) upc_loop_monitor_47;
    upc_loop_intf#(1) upc_loop_intf_48(clock,reset);
    assign upc_loop_intf_48.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_CS_fsm;
    assign upc_loop_intf_48.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_48.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_48.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_48.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_48.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_48.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_48.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_48.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_48.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_48.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_start;
    assign upc_loop_intf_48.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_ready;
    assign upc_loop_intf_48.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_351_1_fu_241.ap_done_int;
    assign upc_loop_intf_48.loop_continue = 1'b1;
    assign upc_loop_intf_48.quit_at_end = 1'b1;
    assign upc_loop_intf_48.finish = finish;
    csv_file_dump upc_loop_csv_dumper_48;
    upc_loop_monitor #(1) upc_loop_monitor_48;
    upc_loop_intf#(1) upc_loop_intf_49(clock,reset);
    assign upc_loop_intf_49.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_CS_fsm;
    assign upc_loop_intf_49.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_49.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_49.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_49.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_49.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_49.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_49.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_49.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_49.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_49.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_start;
    assign upc_loop_intf_49.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_ready;
    assign upc_loop_intf_49.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_1_fu_249.ap_done_int;
    assign upc_loop_intf_49.loop_continue = 1'b1;
    assign upc_loop_intf_49.quit_at_end = 1'b0;
    assign upc_loop_intf_49.finish = finish;
    csv_file_dump upc_loop_csv_dumper_49;
    upc_loop_monitor #(1) upc_loop_monitor_49;
    upc_loop_intf#(1) upc_loop_intf_50(clock,reset);
    assign upc_loop_intf_50.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_CS_fsm;
    assign upc_loop_intf_50.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_50.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_50.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_50.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_50.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_50.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_50.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_50.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_50.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_50.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_start;
    assign upc_loop_intf_50.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_ready;
    assign upc_loop_intf_50.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_360_2_fu_255.ap_done_int;
    assign upc_loop_intf_50.loop_continue = 1'b1;
    assign upc_loop_intf_50.quit_at_end = 1'b0;
    assign upc_loop_intf_50.finish = finish;
    csv_file_dump upc_loop_csv_dumper_50;
    upc_loop_monitor #(1) upc_loop_monitor_50;
    upc_loop_intf#(1) upc_loop_intf_51(clock,reset);
    assign upc_loop_intf_51.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_CS_fsm;
    assign upc_loop_intf_51.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_51.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_51.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_51.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_51.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_51.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_51.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_51.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_51.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_51.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_start;
    assign upc_loop_intf_51.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_ready;
    assign upc_loop_intf_51.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_369_4_fu_273.ap_done_int;
    assign upc_loop_intf_51.loop_continue = 1'b1;
    assign upc_loop_intf_51.quit_at_end = 1'b0;
    assign upc_loop_intf_51.finish = finish;
    csv_file_dump upc_loop_csv_dumper_51;
    upc_loop_monitor #(1) upc_loop_monitor_51;
    upc_loop_intf#(1) upc_loop_intf_52(clock,reset);
    assign upc_loop_intf_52.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_CS_fsm;
    assign upc_loop_intf_52.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_52.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_52.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_52.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_52.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_52.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_52.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_52.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_enable_reg_pp0_iter2;
    assign upc_loop_intf_52.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_52.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_start;
    assign upc_loop_intf_52.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_ready;
    assign upc_loop_intf_52.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_376_5_fu_282.ap_done_int;
    assign upc_loop_intf_52.loop_continue = 1'b1;
    assign upc_loop_intf_52.quit_at_end = 1'b0;
    assign upc_loop_intf_52.finish = finish;
    csv_file_dump upc_loop_csv_dumper_52;
    upc_loop_monitor #(1) upc_loop_monitor_52;
    upc_loop_intf#(1) upc_loop_intf_53(clock,reset);
    assign upc_loop_intf_53.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_CS_fsm;
    assign upc_loop_intf_53.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_53.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_53.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_53.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_53.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_53.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_53.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_53.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_53.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_53.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_start;
    assign upc_loop_intf_53.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_ready;
    assign upc_loop_intf_53.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_shake_absorb_fu_153.grp_shake_absorb_Pipeline_VITIS_LOOP_12_12_fu_308.ap_done_int;
    assign upc_loop_intf_53.loop_continue = 1'b1;
    assign upc_loop_intf_53.quit_at_end = 1'b0;
    assign upc_loop_intf_53.finish = finish;
    csv_file_dump upc_loop_csv_dumper_53;
    upc_loop_monitor #(1) upc_loop_monitor_53;
    upc_loop_intf#(4) upc_loop_intf_54(clock,reset);
    assign upc_loop_intf_54.cur_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_CS_fsm;
    assign upc_loop_intf_54.iter_start_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_54.iter_end_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_54.quit_state = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_54.iter_start_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_54.iter_end_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_54.quit_block = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_54.iter_start_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_54.iter_end_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_54.quit_enable = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_54.loop_start = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_start;
    assign upc_loop_intf_54.loop_ready = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_ready;
    assign upc_loop_intf_54.loop_done = AESL_inst_dpu_keygen.grp_sample_eta_fu_679.grp_sample_eta_Pipeline_VITIS_LOOP_417_2_fu_173.ap_done_int;
    assign upc_loop_intf_54.loop_continue = 1'b1;
    assign upc_loop_intf_54.quit_at_end = 1'b0;
    assign upc_loop_intf_54.finish = finish;
    csv_file_dump upc_loop_csv_dumper_54;
    upc_loop_monitor #(4) upc_loop_monitor_54;
    upc_loop_intf#(1) upc_loop_intf_55(clock,reset);
    assign upc_loop_intf_55.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_CS_fsm;
    assign upc_loop_intf_55.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_55.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_55.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_55.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_55.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_55.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_55.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_55.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_55.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_55.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_start;
    assign upc_loop_intf_55.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_ready;
    assign upc_loop_intf_55.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_17_fu_690.ap_done_int;
    assign upc_loop_intf_55.loop_continue = 1'b1;
    assign upc_loop_intf_55.quit_at_end = 1'b0;
    assign upc_loop_intf_55.finish = finish;
    csv_file_dump upc_loop_csv_dumper_55;
    upc_loop_monitor #(1) upc_loop_monitor_55;
    upc_loop_intf#(1) upc_loop_intf_56(clock,reset);
    assign upc_loop_intf_56.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_CS_fsm;
    assign upc_loop_intf_56.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_56.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_56.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_56.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_56.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_56.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_56.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_56.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_56.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_56.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_start;
    assign upc_loop_intf_56.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_ready;
    assign upc_loop_intf_56.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_18_fu_698.ap_done_int;
    assign upc_loop_intf_56.loop_continue = 1'b1;
    assign upc_loop_intf_56.quit_at_end = 1'b0;
    assign upc_loop_intf_56.finish = finish;
    csv_file_dump upc_loop_csv_dumper_56;
    upc_loop_monitor #(1) upc_loop_monitor_56;
    upc_loop_intf#(1) upc_loop_intf_57(clock,reset);
    assign upc_loop_intf_57.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_CS_fsm;
    assign upc_loop_intf_57.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_57.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_57.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_57.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_57.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_57.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_57.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_57.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_57.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_57.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_start;
    assign upc_loop_intf_57.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_ready;
    assign upc_loop_intf_57.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_55_5_fu_706.ap_done_int;
    assign upc_loop_intf_57.loop_continue = 1'b1;
    assign upc_loop_intf_57.quit_at_end = 1'b0;
    assign upc_loop_intf_57.finish = finish;
    csv_file_dump upc_loop_csv_dumper_57;
    upc_loop_monitor #(1) upc_loop_monitor_57;
    upc_loop_intf#(1) upc_loop_intf_58(clock,reset);
    assign upc_loop_intf_58.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_CS_fsm;
    assign upc_loop_intf_58.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_58.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_58.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_58.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_58.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_58.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_58.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_58.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_58.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_58.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_start;
    assign upc_loop_intf_58.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_ready;
    assign upc_loop_intf_58.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_95_19_fu_719.ap_done_int;
    assign upc_loop_intf_58.loop_continue = 1'b1;
    assign upc_loop_intf_58.quit_at_end = 1'b0;
    assign upc_loop_intf_58.finish = finish;
    csv_file_dump upc_loop_csv_dumper_58;
    upc_loop_monitor #(1) upc_loop_monitor_58;
    upc_loop_intf#(1) upc_loop_intf_59(clock,reset);
    assign upc_loop_intf_59.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_CS_fsm;
    assign upc_loop_intf_59.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_59.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_59.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_59.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_59.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_59.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_59.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_59.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_59.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_59.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_start;
    assign upc_loop_intf_59.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_ready;
    assign upc_loop_intf_59.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_60_6_fu_727.ap_done_int;
    assign upc_loop_intf_59.loop_continue = 1'b1;
    assign upc_loop_intf_59.quit_at_end = 1'b0;
    assign upc_loop_intf_59.finish = finish;
    csv_file_dump upc_loop_csv_dumper_59;
    upc_loop_monitor #(1) upc_loop_monitor_59;
    upc_loop_intf#(1) upc_loop_intf_60(clock,reset);
    assign upc_loop_intf_60.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_CS_fsm;
    assign upc_loop_intf_60.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_60.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_60.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_60.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_60.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_60.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_60.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_60.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_60.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_60.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_start;
    assign upc_loop_intf_60.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_ready;
    assign upc_loop_intf_60.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_61_7_fu_735.ap_done_int;
    assign upc_loop_intf_60.loop_continue = 1'b1;
    assign upc_loop_intf_60.quit_at_end = 1'b0;
    assign upc_loop_intf_60.finish = finish;
    csv_file_dump upc_loop_csv_dumper_60;
    upc_loop_monitor #(1) upc_loop_monitor_60;
    upc_loop_intf#(1) upc_loop_intf_61(clock,reset);
    assign upc_loop_intf_61.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_CS_fsm;
    assign upc_loop_intf_61.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_61.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_61.quit_state = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_61.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_61.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_61.quit_block = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_61.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_61.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_61.quit_enable = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_61.loop_start = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_start;
    assign upc_loop_intf_61.loop_ready = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_ready;
    assign upc_loop_intf_61.loop_done = AESL_inst_dpu_keygen.grp_dpu_pack_fu_743.grp_dpu_pack_Pipeline_VITIS_LOOP_73_1_fu_79.ap_done_int;
    assign upc_loop_intf_61.loop_continue = 1'b1;
    assign upc_loop_intf_61.quit_at_end = 1'b1;
    assign upc_loop_intf_61.finish = finish;
    csv_file_dump upc_loop_csv_dumper_61;
    upc_loop_monitor #(1) upc_loop_monitor_61;
    upc_loop_intf#(4) upc_loop_intf_62(clock,reset);
    assign upc_loop_intf_62.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_CS_fsm;
    assign upc_loop_intf_62.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_62.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_62.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_62.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_62.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_62.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_62.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_62.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_62.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_62.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_start;
    assign upc_loop_intf_62.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_ready;
    assign upc_loop_intf_62.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_369_4_fu_50.ap_done_int;
    assign upc_loop_intf_62.loop_continue = 1'b1;
    assign upc_loop_intf_62.quit_at_end = 1'b0;
    assign upc_loop_intf_62.finish = finish;
    csv_file_dump upc_loop_csv_dumper_62;
    upc_loop_monitor #(4) upc_loop_monitor_62;
    upc_loop_intf#(4) upc_loop_intf_63(clock,reset);
    assign upc_loop_intf_63.cur_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_CS_fsm;
    assign upc_loop_intf_63.iter_start_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_63.iter_end_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_63.quit_state = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_63.iter_start_block = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_63.iter_end_block = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_63.quit_block = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_63.iter_start_enable = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_63.iter_end_enable = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_63.quit_enable = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_63.loop_start = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_start;
    assign upc_loop_intf_63.loop_ready = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_ready;
    assign upc_loop_intf_63.loop_done = AESL_inst_dpu_keygen.grp_shake_absorb_3_fu_752.grp_shake_absorb_3_Pipeline_VITIS_LOOP_376_5_fu_59.ap_done_int;
    assign upc_loop_intf_63.loop_continue = 1'b1;
    assign upc_loop_intf_63.quit_at_end = 1'b0;
    assign upc_loop_intf_63.finish = finish;
    csv_file_dump upc_loop_csv_dumper_63;
    upc_loop_monitor #(4) upc_loop_monitor_63;
    upc_loop_intf#(1) upc_loop_intf_64(clock,reset);
    assign upc_loop_intf_64.cur_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_CS_fsm;
    assign upc_loop_intf_64.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_64.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_64.quit_state = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_64.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_64.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_64.quit_block = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_64.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_64.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_64.quit_enable = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_64.loop_start = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_start;
    assign upc_loop_intf_64.loop_ready = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_ready;
    assign upc_loop_intf_64.loop_done = AESL_inst_dpu_keygen.grp_dpu_keygen_Pipeline_VITIS_LOOP_62_8_fu_769.ap_done_int;
    assign upc_loop_intf_64.loop_continue = 1'b1;
    assign upc_loop_intf_64.quit_at_end = 1'b0;
    assign upc_loop_intf_64.finish = finish;
    csv_file_dump upc_loop_csv_dumper_64;
    upc_loop_monitor #(1) upc_loop_monitor_64;
    upc_loop_intf#(7) upc_loop_intf_65(clock,reset);
    assign upc_loop_intf_65.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_CS_fsm;
    assign upc_loop_intf_65.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_65.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_65.quit_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_ST_fsm_pp0_stage1;
    assign upc_loop_intf_65.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_65.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_65.quit_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_block_pp0_stage1_subdone;
    assign upc_loop_intf_65.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_65.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_65.quit_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_65.loop_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_start;
    assign upc_loop_intf_65.loop_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_ready;
    assign upc_loop_intf_65.loop_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_666_8_fu_234.ap_done_int;
    assign upc_loop_intf_65.loop_continue = 1'b1;
    assign upc_loop_intf_65.quit_at_end = 1'b0;
    assign upc_loop_intf_65.finish = finish;
    csv_file_dump upc_loop_csv_dumper_65;
    upc_loop_monitor #(7) upc_loop_monitor_65;
    upc_loop_intf#(1) upc_loop_intf_66(clock,reset);
    assign upc_loop_intf_66.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_CS_fsm;
    assign upc_loop_intf_66.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_66.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_66.quit_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_66.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_66.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_66.quit_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_66.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_66.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_66.quit_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_66.loop_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_start;
    assign upc_loop_intf_66.loop_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_ready;
    assign upc_loop_intf_66.loop_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_13_fu_252.ap_done_int;
    assign upc_loop_intf_66.loop_continue = 1'b1;
    assign upc_loop_intf_66.quit_at_end = 1'b1;
    assign upc_loop_intf_66.finish = finish;
    csv_file_dump upc_loop_csv_dumper_66;
    upc_loop_monitor #(1) upc_loop_monitor_66;
    upc_loop_intf#(1) upc_loop_intf_67(clock,reset);
    assign upc_loop_intf_67.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_CS_fsm;
    assign upc_loop_intf_67.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_67.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_67.quit_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_67.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_67.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_67.quit_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_67.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_67.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_67.quit_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_67.loop_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_start;
    assign upc_loop_intf_67.loop_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_ready;
    assign upc_loop_intf_67.loop_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_15_fu_269.ap_done_int;
    assign upc_loop_intf_67.loop_continue = 1'b1;
    assign upc_loop_intf_67.quit_at_end = 1'b1;
    assign upc_loop_intf_67.finish = finish;
    csv_file_dump upc_loop_csv_dumper_67;
    upc_loop_monitor #(1) upc_loop_monitor_67;
    upc_loop_intf#(3) upc_loop_intf_68(clock,reset);
    assign upc_loop_intf_68.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_CS_fsm;
    assign upc_loop_intf_68.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_68.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_68.quit_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_68.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_68.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_68.quit_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_68.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_68.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_68.quit_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_68.loop_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_start;
    assign upc_loop_intf_68.loop_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_ready;
    assign upc_loop_intf_68.loop_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_709_12_fu_286.ap_done_int;
    assign upc_loop_intf_68.loop_continue = 1'b1;
    assign upc_loop_intf_68.quit_at_end = 1'b0;
    assign upc_loop_intf_68.finish = finish;
    csv_file_dump upc_loop_csv_dumper_68;
    upc_loop_monitor #(3) upc_loop_monitor_68;
    upc_loop_intf#(1) upc_loop_intf_69(clock,reset);
    assign upc_loop_intf_69.cur_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_CS_fsm;
    assign upc_loop_intf_69.iter_start_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_69.iter_end_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_69.quit_state = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_69.iter_start_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_69.iter_end_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_69.quit_block = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_69.iter_start_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_69.iter_end_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_69.quit_enable = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_enable_reg_pp0_iter1;
    assign upc_loop_intf_69.loop_start = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_start;
    assign upc_loop_intf_69.loop_ready = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_ready;
    assign upc_loop_intf_69.loop_done = AESL_inst_dpu_keygen.grp_dpu_pack_4_fu_776.grp_dpu_pack_4_Pipeline_VITIS_LOOP_73_1_fu_304.ap_done_int;
    assign upc_loop_intf_69.loop_continue = 1'b1;
    assign upc_loop_intf_69.quit_at_end = 1'b1;
    assign upc_loop_intf_69.finish = finish;
    csv_file_dump upc_loop_csv_dumper_69;
    upc_loop_monitor #(1) upc_loop_monitor_69;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);
    mstatus_csv_dumper_53 = new("./module_status53.csv");
    module_monitor_53 = new(module_intf_53,mstatus_csv_dumper_53);
    mstatus_csv_dumper_54 = new("./module_status54.csv");
    module_monitor_54 = new(module_intf_54,mstatus_csv_dumper_54);
    mstatus_csv_dumper_55 = new("./module_status55.csv");
    module_monitor_55 = new(module_intf_55,mstatus_csv_dumper_55);
    mstatus_csv_dumper_56 = new("./module_status56.csv");
    module_monitor_56 = new(module_intf_56,mstatus_csv_dumper_56);
    mstatus_csv_dumper_57 = new("./module_status57.csv");
    module_monitor_57 = new(module_intf_57,mstatus_csv_dumper_57);
    mstatus_csv_dumper_58 = new("./module_status58.csv");
    module_monitor_58 = new(module_intf_58,mstatus_csv_dumper_58);
    mstatus_csv_dumper_59 = new("./module_status59.csv");
    module_monitor_59 = new(module_intf_59,mstatus_csv_dumper_59);
    mstatus_csv_dumper_60 = new("./module_status60.csv");
    module_monitor_60 = new(module_intf_60,mstatus_csv_dumper_60);
    mstatus_csv_dumper_61 = new("./module_status61.csv");
    module_monitor_61 = new(module_intf_61,mstatus_csv_dumper_61);
    mstatus_csv_dumper_62 = new("./module_status62.csv");
    module_monitor_62 = new(module_intf_62,mstatus_csv_dumper_62);
    mstatus_csv_dumper_63 = new("./module_status63.csv");
    module_monitor_63 = new(module_intf_63,mstatus_csv_dumper_63);
    mstatus_csv_dumper_64 = new("./module_status64.csv");
    module_monitor_64 = new(module_intf_64,mstatus_csv_dumper_64);
    mstatus_csv_dumper_65 = new("./module_status65.csv");
    module_monitor_65 = new(module_intf_65,mstatus_csv_dumper_65);
    mstatus_csv_dumper_66 = new("./module_status66.csv");
    module_monitor_66 = new(module_intf_66,mstatus_csv_dumper_66);
    mstatus_csv_dumper_67 = new("./module_status67.csv");
    module_monitor_67 = new(module_intf_67,mstatus_csv_dumper_67);
    mstatus_csv_dumper_68 = new("./module_status68.csv");
    module_monitor_68 = new(module_intf_68,mstatus_csv_dumper_68);
    mstatus_csv_dumper_69 = new("./module_status69.csv");
    module_monitor_69 = new(module_intf_69,mstatus_csv_dumper_69);
    mstatus_csv_dumper_70 = new("./module_status70.csv");
    module_monitor_70 = new(module_intf_70,mstatus_csv_dumper_70);
    mstatus_csv_dumper_71 = new("./module_status71.csv");
    module_monitor_71 = new(module_intf_71,mstatus_csv_dumper_71);
    mstatus_csv_dumper_72 = new("./module_status72.csv");
    module_monitor_72 = new(module_intf_72,mstatus_csv_dumper_72);
    mstatus_csv_dumper_73 = new("./module_status73.csv");
    module_monitor_73 = new(module_intf_73,mstatus_csv_dumper_73);
    mstatus_csv_dumper_74 = new("./module_status74.csv");
    module_monitor_74 = new(module_intf_74,mstatus_csv_dumper_74);
    mstatus_csv_dumper_75 = new("./module_status75.csv");
    module_monitor_75 = new(module_intf_75,mstatus_csv_dumper_75);
    mstatus_csv_dumper_76 = new("./module_status76.csv");
    module_monitor_76 = new(module_intf_76,mstatus_csv_dumper_76);
    mstatus_csv_dumper_77 = new("./module_status77.csv");
    module_monitor_77 = new(module_intf_77,mstatus_csv_dumper_77);
    mstatus_csv_dumper_78 = new("./module_status78.csv");
    module_monitor_78 = new(module_intf_78,mstatus_csv_dumper_78);
    mstatus_csv_dumper_79 = new("./module_status79.csv");
    module_monitor_79 = new(module_intf_79,mstatus_csv_dumper_79);
    mstatus_csv_dumper_80 = new("./module_status80.csv");
    module_monitor_80 = new(module_intf_80,mstatus_csv_dumper_80);
    mstatus_csv_dumper_81 = new("./module_status81.csv");
    module_monitor_81 = new(module_intf_81,mstatus_csv_dumper_81);
    mstatus_csv_dumper_82 = new("./module_status82.csv");
    module_monitor_82 = new(module_intf_82,mstatus_csv_dumper_82);
    mstatus_csv_dumper_83 = new("./module_status83.csv");
    module_monitor_83 = new(module_intf_83,mstatus_csv_dumper_83);
    mstatus_csv_dumper_84 = new("./module_status84.csv");
    module_monitor_84 = new(module_intf_84,mstatus_csv_dumper_84);
    mstatus_csv_dumper_85 = new("./module_status85.csv");
    module_monitor_85 = new(module_intf_85,mstatus_csv_dumper_85);
    mstatus_csv_dumper_86 = new("./module_status86.csv");
    module_monitor_86 = new(module_intf_86,mstatus_csv_dumper_86);
    mstatus_csv_dumper_87 = new("./module_status87.csv");
    module_monitor_87 = new(module_intf_87,mstatus_csv_dumper_87);
    mstatus_csv_dumper_88 = new("./module_status88.csv");
    module_monitor_88 = new(module_intf_88,mstatus_csv_dumper_88);
    mstatus_csv_dumper_89 = new("./module_status89.csv");
    module_monitor_89 = new(module_intf_89,mstatus_csv_dumper_89);
    mstatus_csv_dumper_90 = new("./module_status90.csv");
    module_monitor_90 = new(module_intf_90,mstatus_csv_dumper_90);
    mstatus_csv_dumper_91 = new("./module_status91.csv");
    module_monitor_91 = new(module_intf_91,mstatus_csv_dumper_91);
    mstatus_csv_dumper_92 = new("./module_status92.csv");
    module_monitor_92 = new(module_intf_92,mstatus_csv_dumper_92);
    mstatus_csv_dumper_93 = new("./module_status93.csv");
    module_monitor_93 = new(module_intf_93,mstatus_csv_dumper_93);
    mstatus_csv_dumper_94 = new("./module_status94.csv");
    module_monitor_94 = new(module_intf_94,mstatus_csv_dumper_94);
    mstatus_csv_dumper_95 = new("./module_status95.csv");
    module_monitor_95 = new(module_intf_95,mstatus_csv_dumper_95);
    mstatus_csv_dumper_96 = new("./module_status96.csv");
    module_monitor_96 = new(module_intf_96,mstatus_csv_dumper_96);
    mstatus_csv_dumper_97 = new("./module_status97.csv");
    module_monitor_97 = new(module_intf_97,mstatus_csv_dumper_97);
    mstatus_csv_dumper_98 = new("./module_status98.csv");
    module_monitor_98 = new(module_intf_98,mstatus_csv_dumper_98);
    mstatus_csv_dumper_99 = new("./module_status99.csv");
    module_monitor_99 = new(module_intf_99,mstatus_csv_dumper_99);
    mstatus_csv_dumper_100 = new("./module_status100.csv");
    module_monitor_100 = new(module_intf_100,mstatus_csv_dumper_100);
    mstatus_csv_dumper_101 = new("./module_status101.csv");
    module_monitor_101 = new(module_intf_101,mstatus_csv_dumper_101);
    mstatus_csv_dumper_102 = new("./module_status102.csv");
    module_monitor_102 = new(module_intf_102,mstatus_csv_dumper_102);
    mstatus_csv_dumper_103 = new("./module_status103.csv");
    module_monitor_103 = new(module_intf_103,mstatus_csv_dumper_103);
    mstatus_csv_dumper_104 = new("./module_status104.csv");
    module_monitor_104 = new(module_intf_104,mstatus_csv_dumper_104);
    mstatus_csv_dumper_105 = new("./module_status105.csv");
    module_monitor_105 = new(module_intf_105,mstatus_csv_dumper_105);
    mstatus_csv_dumper_106 = new("./module_status106.csv");
    module_monitor_106 = new(module_intf_106,mstatus_csv_dumper_106);
    mstatus_csv_dumper_107 = new("./module_status107.csv");
    module_monitor_107 = new(module_intf_107,mstatus_csv_dumper_107);
    mstatus_csv_dumper_108 = new("./module_status108.csv");
    module_monitor_108 = new(module_intf_108,mstatus_csv_dumper_108);
    mstatus_csv_dumper_109 = new("./module_status109.csv");
    module_monitor_109 = new(module_intf_109,mstatus_csv_dumper_109);
    mstatus_csv_dumper_110 = new("./module_status110.csv");
    module_monitor_110 = new(module_intf_110,mstatus_csv_dumper_110);
    mstatus_csv_dumper_111 = new("./module_status111.csv");
    module_monitor_111 = new(module_intf_111,mstatus_csv_dumper_111);
    mstatus_csv_dumper_112 = new("./module_status112.csv");
    module_monitor_112 = new(module_intf_112,mstatus_csv_dumper_112);
    mstatus_csv_dumper_113 = new("./module_status113.csv");
    module_monitor_113 = new(module_intf_113,mstatus_csv_dumper_113);
    mstatus_csv_dumper_114 = new("./module_status114.csv");
    module_monitor_114 = new(module_intf_114,mstatus_csv_dumper_114);
    mstatus_csv_dumper_115 = new("./module_status115.csv");
    module_monitor_115 = new(module_intf_115,mstatus_csv_dumper_115);
    mstatus_csv_dumper_116 = new("./module_status116.csv");
    module_monitor_116 = new(module_intf_116,mstatus_csv_dumper_116);
    mstatus_csv_dumper_117 = new("./module_status117.csv");
    module_monitor_117 = new(module_intf_117,mstatus_csv_dumper_117);
    mstatus_csv_dumper_118 = new("./module_status118.csv");
    module_monitor_118 = new(module_intf_118,mstatus_csv_dumper_118);
    mstatus_csv_dumper_119 = new("./module_status119.csv");
    module_monitor_119 = new(module_intf_119,mstatus_csv_dumper_119);
    mstatus_csv_dumper_120 = new("./module_status120.csv");
    module_monitor_120 = new(module_intf_120,mstatus_csv_dumper_120);
    mstatus_csv_dumper_121 = new("./module_status121.csv");
    module_monitor_121 = new(module_intf_121,mstatus_csv_dumper_121);
    mstatus_csv_dumper_122 = new("./module_status122.csv");
    module_monitor_122 = new(module_intf_122,mstatus_csv_dumper_122);
    mstatus_csv_dumper_123 = new("./module_status123.csv");
    module_monitor_123 = new(module_intf_123,mstatus_csv_dumper_123);
    mstatus_csv_dumper_124 = new("./module_status124.csv");
    module_monitor_124 = new(module_intf_124,mstatus_csv_dumper_124);
    mstatus_csv_dumper_125 = new("./module_status125.csv");
    module_monitor_125 = new(module_intf_125,mstatus_csv_dumper_125);
    mstatus_csv_dumper_126 = new("./module_status126.csv");
    module_monitor_126 = new(module_intf_126,mstatus_csv_dumper_126);
    mstatus_csv_dumper_127 = new("./module_status127.csv");
    module_monitor_127 = new(module_intf_127,mstatus_csv_dumper_127);
    mstatus_csv_dumper_128 = new("./module_status128.csv");
    module_monitor_128 = new(module_intf_128,mstatus_csv_dumper_128);
    mstatus_csv_dumper_129 = new("./module_status129.csv");
    module_monitor_129 = new(module_intf_129,mstatus_csv_dumper_129);
    mstatus_csv_dumper_130 = new("./module_status130.csv");
    module_monitor_130 = new(module_intf_130,mstatus_csv_dumper_130);
    mstatus_csv_dumper_131 = new("./module_status131.csv");
    module_monitor_131 = new(module_intf_131,mstatus_csv_dumper_131);
    mstatus_csv_dumper_132 = new("./module_status132.csv");
    module_monitor_132 = new(module_intf_132,mstatus_csv_dumper_132);
    mstatus_csv_dumper_133 = new("./module_status133.csv");
    module_monitor_133 = new(module_intf_133,mstatus_csv_dumper_133);
    mstatus_csv_dumper_134 = new("./module_status134.csv");
    module_monitor_134 = new(module_intf_134,mstatus_csv_dumper_134);
    mstatus_csv_dumper_135 = new("./module_status135.csv");
    module_monitor_135 = new(module_intf_135,mstatus_csv_dumper_135);
    mstatus_csv_dumper_136 = new("./module_status136.csv");
    module_monitor_136 = new(module_intf_136,mstatus_csv_dumper_136);
    mstatus_csv_dumper_137 = new("./module_status137.csv");
    module_monitor_137 = new(module_intf_137,mstatus_csv_dumper_137);
    mstatus_csv_dumper_138 = new("./module_status138.csv");
    module_monitor_138 = new(module_intf_138,mstatus_csv_dumper_138);
    mstatus_csv_dumper_139 = new("./module_status139.csv");
    module_monitor_139 = new(module_intf_139,mstatus_csv_dumper_139);
    mstatus_csv_dumper_140 = new("./module_status140.csv");
    module_monitor_140 = new(module_intf_140,mstatus_csv_dumper_140);
    mstatus_csv_dumper_141 = new("./module_status141.csv");
    module_monitor_141 = new(module_intf_141,mstatus_csv_dumper_141);
    mstatus_csv_dumper_142 = new("./module_status142.csv");
    module_monitor_142 = new(module_intf_142,mstatus_csv_dumper_142);
    mstatus_csv_dumper_143 = new("./module_status143.csv");
    module_monitor_143 = new(module_intf_143,mstatus_csv_dumper_143);
    mstatus_csv_dumper_144 = new("./module_status144.csv");
    module_monitor_144 = new(module_intf_144,mstatus_csv_dumper_144);
    mstatus_csv_dumper_145 = new("./module_status145.csv");
    module_monitor_145 = new(module_intf_145,mstatus_csv_dumper_145);
    mstatus_csv_dumper_146 = new("./module_status146.csv");
    module_monitor_146 = new(module_intf_146,mstatus_csv_dumper_146);
    mstatus_csv_dumper_147 = new("./module_status147.csv");
    module_monitor_147 = new(module_intf_147,mstatus_csv_dumper_147);
    mstatus_csv_dumper_148 = new("./module_status148.csv");
    module_monitor_148 = new(module_intf_148,mstatus_csv_dumper_148);
    mstatus_csv_dumper_149 = new("./module_status149.csv");
    module_monitor_149 = new(module_intf_149,mstatus_csv_dumper_149);
    mstatus_csv_dumper_150 = new("./module_status150.csv");
    module_monitor_150 = new(module_intf_150,mstatus_csv_dumper_150);
    mstatus_csv_dumper_151 = new("./module_status151.csv");
    module_monitor_151 = new(module_intf_151,mstatus_csv_dumper_151);
    mstatus_csv_dumper_152 = new("./module_status152.csv");
    module_monitor_152 = new(module_intf_152,mstatus_csv_dumper_152);
    mstatus_csv_dumper_153 = new("./module_status153.csv");
    module_monitor_153 = new(module_intf_153,mstatus_csv_dumper_153);
    mstatus_csv_dumper_154 = new("./module_status154.csv");
    module_monitor_154 = new(module_intf_154,mstatus_csv_dumper_154);
    mstatus_csv_dumper_155 = new("./module_status155.csv");
    module_monitor_155 = new(module_intf_155,mstatus_csv_dumper_155);
    mstatus_csv_dumper_156 = new("./module_status156.csv");
    module_monitor_156 = new(module_intf_156,mstatus_csv_dumper_156);
    mstatus_csv_dumper_157 = new("./module_status157.csv");
    module_monitor_157 = new(module_intf_157,mstatus_csv_dumper_157);
    mstatus_csv_dumper_158 = new("./module_status158.csv");
    module_monitor_158 = new(module_intf_158,mstatus_csv_dumper_158);
    mstatus_csv_dumper_159 = new("./module_status159.csv");
    module_monitor_159 = new(module_intf_159,mstatus_csv_dumper_159);
    mstatus_csv_dumper_160 = new("./module_status160.csv");
    module_monitor_160 = new(module_intf_160,mstatus_csv_dumper_160);
    mstatus_csv_dumper_161 = new("./module_status161.csv");
    module_monitor_161 = new(module_intf_161,mstatus_csv_dumper_161);
    mstatus_csv_dumper_162 = new("./module_status162.csv");
    module_monitor_162 = new(module_intf_162,mstatus_csv_dumper_162);
    mstatus_csv_dumper_163 = new("./module_status163.csv");
    module_monitor_163 = new(module_intf_163,mstatus_csv_dumper_163);
    mstatus_csv_dumper_164 = new("./module_status164.csv");
    module_monitor_164 = new(module_intf_164,mstatus_csv_dumper_164);
    mstatus_csv_dumper_165 = new("./module_status165.csv");
    module_monitor_165 = new(module_intf_165,mstatus_csv_dumper_165);
    mstatus_csv_dumper_166 = new("./module_status166.csv");
    module_monitor_166 = new(module_intf_166,mstatus_csv_dumper_166);
    mstatus_csv_dumper_167 = new("./module_status167.csv");
    module_monitor_167 = new(module_intf_167,mstatus_csv_dumper_167);
    mstatus_csv_dumper_168 = new("./module_status168.csv");
    module_monitor_168 = new(module_intf_168,mstatus_csv_dumper_168);
    mstatus_csv_dumper_169 = new("./module_status169.csv");
    module_monitor_169 = new(module_intf_169,mstatus_csv_dumper_169);
    mstatus_csv_dumper_170 = new("./module_status170.csv");
    module_monitor_170 = new(module_intf_170,mstatus_csv_dumper_170);
    mstatus_csv_dumper_171 = new("./module_status171.csv");
    module_monitor_171 = new(module_intf_171,mstatus_csv_dumper_171);
    mstatus_csv_dumper_172 = new("./module_status172.csv");
    module_monitor_172 = new(module_intf_172,mstatus_csv_dumper_172);
    mstatus_csv_dumper_173 = new("./module_status173.csv");
    module_monitor_173 = new(module_intf_173,mstatus_csv_dumper_173);
    mstatus_csv_dumper_174 = new("./module_status174.csv");
    module_monitor_174 = new(module_intf_174,mstatus_csv_dumper_174);
    mstatus_csv_dumper_175 = new("./module_status175.csv");
    module_monitor_175 = new(module_intf_175,mstatus_csv_dumper_175);
    mstatus_csv_dumper_176 = new("./module_status176.csv");
    module_monitor_176 = new(module_intf_176,mstatus_csv_dumper_176);
    mstatus_csv_dumper_177 = new("./module_status177.csv");
    module_monitor_177 = new(module_intf_177,mstatus_csv_dumper_177);
    mstatus_csv_dumper_178 = new("./module_status178.csv");
    module_monitor_178 = new(module_intf_178,mstatus_csv_dumper_178);
    mstatus_csv_dumper_179 = new("./module_status179.csv");
    module_monitor_179 = new(module_intf_179,mstatus_csv_dumper_179);
    mstatus_csv_dumper_180 = new("./module_status180.csv");
    module_monitor_180 = new(module_intf_180,mstatus_csv_dumper_180);

    pp_loop_csv_dumper_1 = new("./pp_loop_status1.csv");
    pp_loop_monitor_1 = new(pp_loop_intf_1,pp_loop_csv_dumper_1);
    pp_loop_csv_dumper_2 = new("./pp_loop_status2.csv");
    pp_loop_monitor_2 = new(pp_loop_intf_2,pp_loop_csv_dumper_2);
    pp_loop_csv_dumper_3 = new("./pp_loop_status3.csv");
    pp_loop_monitor_3 = new(pp_loop_intf_3,pp_loop_csv_dumper_3);


    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);
    seq_loop_csv_dumper_10 = new("./seq_loop_status10.csv");
    seq_loop_monitor_10 = new(seq_loop_intf_10,seq_loop_csv_dumper_10);
    seq_loop_csv_dumper_11 = new("./seq_loop_status11.csv");
    seq_loop_monitor_11 = new(seq_loop_intf_11,seq_loop_csv_dumper_11);
    seq_loop_csv_dumper_12 = new("./seq_loop_status12.csv");
    seq_loop_monitor_12 = new(seq_loop_intf_12,seq_loop_csv_dumper_12);
    seq_loop_csv_dumper_13 = new("./seq_loop_status13.csv");
    seq_loop_monitor_13 = new(seq_loop_intf_13,seq_loop_csv_dumper_13);
    seq_loop_csv_dumper_14 = new("./seq_loop_status14.csv");
    seq_loop_monitor_14 = new(seq_loop_intf_14,seq_loop_csv_dumper_14);
    seq_loop_csv_dumper_15 = new("./seq_loop_status15.csv");
    seq_loop_monitor_15 = new(seq_loop_intf_15,seq_loop_csv_dumper_15);
    seq_loop_csv_dumper_16 = new("./seq_loop_status16.csv");
    seq_loop_monitor_16 = new(seq_loop_intf_16,seq_loop_csv_dumper_16);
    seq_loop_csv_dumper_17 = new("./seq_loop_status17.csv");
    seq_loop_monitor_17 = new(seq_loop_intf_17,seq_loop_csv_dumper_17);
    seq_loop_csv_dumper_18 = new("./seq_loop_status18.csv");
    seq_loop_monitor_18 = new(seq_loop_intf_18,seq_loop_csv_dumper_18);
    seq_loop_csv_dumper_19 = new("./seq_loop_status19.csv");
    seq_loop_monitor_19 = new(seq_loop_intf_19,seq_loop_csv_dumper_19);
    seq_loop_csv_dumper_20 = new("./seq_loop_status20.csv");
    seq_loop_monitor_20 = new(seq_loop_intf_20,seq_loop_csv_dumper_20);
    seq_loop_csv_dumper_21 = new("./seq_loop_status21.csv");
    seq_loop_monitor_21 = new(seq_loop_intf_21,seq_loop_csv_dumper_21);
    seq_loop_csv_dumper_22 = new("./seq_loop_status22.csv");
    seq_loop_monitor_22 = new(seq_loop_intf_22,seq_loop_csv_dumper_22);
    seq_loop_csv_dumper_23 = new("./seq_loop_status23.csv");
    seq_loop_monitor_23 = new(seq_loop_intf_23,seq_loop_csv_dumper_23);
    seq_loop_csv_dumper_24 = new("./seq_loop_status24.csv");
    seq_loop_monitor_24 = new(seq_loop_intf_24,seq_loop_csv_dumper_24);
    seq_loop_csv_dumper_25 = new("./seq_loop_status25.csv");
    seq_loop_monitor_25 = new(seq_loop_intf_25,seq_loop_csv_dumper_25);
    seq_loop_csv_dumper_26 = new("./seq_loop_status26.csv");
    seq_loop_monitor_26 = new(seq_loop_intf_26,seq_loop_csv_dumper_26);
    seq_loop_csv_dumper_27 = new("./seq_loop_status27.csv");
    seq_loop_monitor_27 = new(seq_loop_intf_27,seq_loop_csv_dumper_27);
    seq_loop_csv_dumper_28 = new("./seq_loop_status28.csv");
    seq_loop_monitor_28 = new(seq_loop_intf_28,seq_loop_csv_dumper_28);
    seq_loop_csv_dumper_29 = new("./seq_loop_status29.csv");
    seq_loop_monitor_29 = new(seq_loop_intf_29,seq_loop_csv_dumper_29);
    seq_loop_csv_dumper_30 = new("./seq_loop_status30.csv");
    seq_loop_monitor_30 = new(seq_loop_intf_30,seq_loop_csv_dumper_30);
    seq_loop_csv_dumper_31 = new("./seq_loop_status31.csv");
    seq_loop_monitor_31 = new(seq_loop_intf_31,seq_loop_csv_dumper_31);
    seq_loop_csv_dumper_32 = new("./seq_loop_status32.csv");
    seq_loop_monitor_32 = new(seq_loop_intf_32,seq_loop_csv_dumper_32);
    seq_loop_csv_dumper_33 = new("./seq_loop_status33.csv");
    seq_loop_monitor_33 = new(seq_loop_intf_33,seq_loop_csv_dumper_33);
    seq_loop_csv_dumper_34 = new("./seq_loop_status34.csv");
    seq_loop_monitor_34 = new(seq_loop_intf_34,seq_loop_csv_dumper_34);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);
    upc_loop_csv_dumper_2 = new("./upc_loop_status2.csv");
    upc_loop_monitor_2 = new(upc_loop_intf_2,upc_loop_csv_dumper_2);
    upc_loop_csv_dumper_3 = new("./upc_loop_status3.csv");
    upc_loop_monitor_3 = new(upc_loop_intf_3,upc_loop_csv_dumper_3);
    upc_loop_csv_dumper_4 = new("./upc_loop_status4.csv");
    upc_loop_monitor_4 = new(upc_loop_intf_4,upc_loop_csv_dumper_4);
    upc_loop_csv_dumper_5 = new("./upc_loop_status5.csv");
    upc_loop_monitor_5 = new(upc_loop_intf_5,upc_loop_csv_dumper_5);
    upc_loop_csv_dumper_6 = new("./upc_loop_status6.csv");
    upc_loop_monitor_6 = new(upc_loop_intf_6,upc_loop_csv_dumper_6);
    upc_loop_csv_dumper_7 = new("./upc_loop_status7.csv");
    upc_loop_monitor_7 = new(upc_loop_intf_7,upc_loop_csv_dumper_7);
    upc_loop_csv_dumper_8 = new("./upc_loop_status8.csv");
    upc_loop_monitor_8 = new(upc_loop_intf_8,upc_loop_csv_dumper_8);
    upc_loop_csv_dumper_9 = new("./upc_loop_status9.csv");
    upc_loop_monitor_9 = new(upc_loop_intf_9,upc_loop_csv_dumper_9);
    upc_loop_csv_dumper_10 = new("./upc_loop_status10.csv");
    upc_loop_monitor_10 = new(upc_loop_intf_10,upc_loop_csv_dumper_10);
    upc_loop_csv_dumper_11 = new("./upc_loop_status11.csv");
    upc_loop_monitor_11 = new(upc_loop_intf_11,upc_loop_csv_dumper_11);
    upc_loop_csv_dumper_12 = new("./upc_loop_status12.csv");
    upc_loop_monitor_12 = new(upc_loop_intf_12,upc_loop_csv_dumper_12);
    upc_loop_csv_dumper_13 = new("./upc_loop_status13.csv");
    upc_loop_monitor_13 = new(upc_loop_intf_13,upc_loop_csv_dumper_13);
    upc_loop_csv_dumper_14 = new("./upc_loop_status14.csv");
    upc_loop_monitor_14 = new(upc_loop_intf_14,upc_loop_csv_dumper_14);
    upc_loop_csv_dumper_15 = new("./upc_loop_status15.csv");
    upc_loop_monitor_15 = new(upc_loop_intf_15,upc_loop_csv_dumper_15);
    upc_loop_csv_dumper_16 = new("./upc_loop_status16.csv");
    upc_loop_monitor_16 = new(upc_loop_intf_16,upc_loop_csv_dumper_16);
    upc_loop_csv_dumper_17 = new("./upc_loop_status17.csv");
    upc_loop_monitor_17 = new(upc_loop_intf_17,upc_loop_csv_dumper_17);
    upc_loop_csv_dumper_18 = new("./upc_loop_status18.csv");
    upc_loop_monitor_18 = new(upc_loop_intf_18,upc_loop_csv_dumper_18);
    upc_loop_csv_dumper_19 = new("./upc_loop_status19.csv");
    upc_loop_monitor_19 = new(upc_loop_intf_19,upc_loop_csv_dumper_19);
    upc_loop_csv_dumper_20 = new("./upc_loop_status20.csv");
    upc_loop_monitor_20 = new(upc_loop_intf_20,upc_loop_csv_dumper_20);
    upc_loop_csv_dumper_21 = new("./upc_loop_status21.csv");
    upc_loop_monitor_21 = new(upc_loop_intf_21,upc_loop_csv_dumper_21);
    upc_loop_csv_dumper_22 = new("./upc_loop_status22.csv");
    upc_loop_monitor_22 = new(upc_loop_intf_22,upc_loop_csv_dumper_22);
    upc_loop_csv_dumper_23 = new("./upc_loop_status23.csv");
    upc_loop_monitor_23 = new(upc_loop_intf_23,upc_loop_csv_dumper_23);
    upc_loop_csv_dumper_24 = new("./upc_loop_status24.csv");
    upc_loop_monitor_24 = new(upc_loop_intf_24,upc_loop_csv_dumper_24);
    upc_loop_csv_dumper_25 = new("./upc_loop_status25.csv");
    upc_loop_monitor_25 = new(upc_loop_intf_25,upc_loop_csv_dumper_25);
    upc_loop_csv_dumper_26 = new("./upc_loop_status26.csv");
    upc_loop_monitor_26 = new(upc_loop_intf_26,upc_loop_csv_dumper_26);
    upc_loop_csv_dumper_27 = new("./upc_loop_status27.csv");
    upc_loop_monitor_27 = new(upc_loop_intf_27,upc_loop_csv_dumper_27);
    upc_loop_csv_dumper_28 = new("./upc_loop_status28.csv");
    upc_loop_monitor_28 = new(upc_loop_intf_28,upc_loop_csv_dumper_28);
    upc_loop_csv_dumper_29 = new("./upc_loop_status29.csv");
    upc_loop_monitor_29 = new(upc_loop_intf_29,upc_loop_csv_dumper_29);
    upc_loop_csv_dumper_30 = new("./upc_loop_status30.csv");
    upc_loop_monitor_30 = new(upc_loop_intf_30,upc_loop_csv_dumper_30);
    upc_loop_csv_dumper_31 = new("./upc_loop_status31.csv");
    upc_loop_monitor_31 = new(upc_loop_intf_31,upc_loop_csv_dumper_31);
    upc_loop_csv_dumper_32 = new("./upc_loop_status32.csv");
    upc_loop_monitor_32 = new(upc_loop_intf_32,upc_loop_csv_dumper_32);
    upc_loop_csv_dumper_33 = new("./upc_loop_status33.csv");
    upc_loop_monitor_33 = new(upc_loop_intf_33,upc_loop_csv_dumper_33);
    upc_loop_csv_dumper_34 = new("./upc_loop_status34.csv");
    upc_loop_monitor_34 = new(upc_loop_intf_34,upc_loop_csv_dumper_34);
    upc_loop_csv_dumper_35 = new("./upc_loop_status35.csv");
    upc_loop_monitor_35 = new(upc_loop_intf_35,upc_loop_csv_dumper_35);
    upc_loop_csv_dumper_36 = new("./upc_loop_status36.csv");
    upc_loop_monitor_36 = new(upc_loop_intf_36,upc_loop_csv_dumper_36);
    upc_loop_csv_dumper_37 = new("./upc_loop_status37.csv");
    upc_loop_monitor_37 = new(upc_loop_intf_37,upc_loop_csv_dumper_37);
    upc_loop_csv_dumper_38 = new("./upc_loop_status38.csv");
    upc_loop_monitor_38 = new(upc_loop_intf_38,upc_loop_csv_dumper_38);
    upc_loop_csv_dumper_39 = new("./upc_loop_status39.csv");
    upc_loop_monitor_39 = new(upc_loop_intf_39,upc_loop_csv_dumper_39);
    upc_loop_csv_dumper_40 = new("./upc_loop_status40.csv");
    upc_loop_monitor_40 = new(upc_loop_intf_40,upc_loop_csv_dumper_40);
    upc_loop_csv_dumper_41 = new("./upc_loop_status41.csv");
    upc_loop_monitor_41 = new(upc_loop_intf_41,upc_loop_csv_dumper_41);
    upc_loop_csv_dumper_42 = new("./upc_loop_status42.csv");
    upc_loop_monitor_42 = new(upc_loop_intf_42,upc_loop_csv_dumper_42);
    upc_loop_csv_dumper_43 = new("./upc_loop_status43.csv");
    upc_loop_monitor_43 = new(upc_loop_intf_43,upc_loop_csv_dumper_43);
    upc_loop_csv_dumper_44 = new("./upc_loop_status44.csv");
    upc_loop_monitor_44 = new(upc_loop_intf_44,upc_loop_csv_dumper_44);
    upc_loop_csv_dumper_45 = new("./upc_loop_status45.csv");
    upc_loop_monitor_45 = new(upc_loop_intf_45,upc_loop_csv_dumper_45);
    upc_loop_csv_dumper_46 = new("./upc_loop_status46.csv");
    upc_loop_monitor_46 = new(upc_loop_intf_46,upc_loop_csv_dumper_46);
    upc_loop_csv_dumper_47 = new("./upc_loop_status47.csv");
    upc_loop_monitor_47 = new(upc_loop_intf_47,upc_loop_csv_dumper_47);
    upc_loop_csv_dumper_48 = new("./upc_loop_status48.csv");
    upc_loop_monitor_48 = new(upc_loop_intf_48,upc_loop_csv_dumper_48);
    upc_loop_csv_dumper_49 = new("./upc_loop_status49.csv");
    upc_loop_monitor_49 = new(upc_loop_intf_49,upc_loop_csv_dumper_49);
    upc_loop_csv_dumper_50 = new("./upc_loop_status50.csv");
    upc_loop_monitor_50 = new(upc_loop_intf_50,upc_loop_csv_dumper_50);
    upc_loop_csv_dumper_51 = new("./upc_loop_status51.csv");
    upc_loop_monitor_51 = new(upc_loop_intf_51,upc_loop_csv_dumper_51);
    upc_loop_csv_dumper_52 = new("./upc_loop_status52.csv");
    upc_loop_monitor_52 = new(upc_loop_intf_52,upc_loop_csv_dumper_52);
    upc_loop_csv_dumper_53 = new("./upc_loop_status53.csv");
    upc_loop_monitor_53 = new(upc_loop_intf_53,upc_loop_csv_dumper_53);
    upc_loop_csv_dumper_54 = new("./upc_loop_status54.csv");
    upc_loop_monitor_54 = new(upc_loop_intf_54,upc_loop_csv_dumper_54);
    upc_loop_csv_dumper_55 = new("./upc_loop_status55.csv");
    upc_loop_monitor_55 = new(upc_loop_intf_55,upc_loop_csv_dumper_55);
    upc_loop_csv_dumper_56 = new("./upc_loop_status56.csv");
    upc_loop_monitor_56 = new(upc_loop_intf_56,upc_loop_csv_dumper_56);
    upc_loop_csv_dumper_57 = new("./upc_loop_status57.csv");
    upc_loop_monitor_57 = new(upc_loop_intf_57,upc_loop_csv_dumper_57);
    upc_loop_csv_dumper_58 = new("./upc_loop_status58.csv");
    upc_loop_monitor_58 = new(upc_loop_intf_58,upc_loop_csv_dumper_58);
    upc_loop_csv_dumper_59 = new("./upc_loop_status59.csv");
    upc_loop_monitor_59 = new(upc_loop_intf_59,upc_loop_csv_dumper_59);
    upc_loop_csv_dumper_60 = new("./upc_loop_status60.csv");
    upc_loop_monitor_60 = new(upc_loop_intf_60,upc_loop_csv_dumper_60);
    upc_loop_csv_dumper_61 = new("./upc_loop_status61.csv");
    upc_loop_monitor_61 = new(upc_loop_intf_61,upc_loop_csv_dumper_61);
    upc_loop_csv_dumper_62 = new("./upc_loop_status62.csv");
    upc_loop_monitor_62 = new(upc_loop_intf_62,upc_loop_csv_dumper_62);
    upc_loop_csv_dumper_63 = new("./upc_loop_status63.csv");
    upc_loop_monitor_63 = new(upc_loop_intf_63,upc_loop_csv_dumper_63);
    upc_loop_csv_dumper_64 = new("./upc_loop_status64.csv");
    upc_loop_monitor_64 = new(upc_loop_intf_64,upc_loop_csv_dumper_64);
    upc_loop_csv_dumper_65 = new("./upc_loop_status65.csv");
    upc_loop_monitor_65 = new(upc_loop_intf_65,upc_loop_csv_dumper_65);
    upc_loop_csv_dumper_66 = new("./upc_loop_status66.csv");
    upc_loop_monitor_66 = new(upc_loop_intf_66,upc_loop_csv_dumper_66);
    upc_loop_csv_dumper_67 = new("./upc_loop_status67.csv");
    upc_loop_monitor_67 = new(upc_loop_intf_67,upc_loop_csv_dumper_67);
    upc_loop_csv_dumper_68 = new("./upc_loop_status68.csv");
    upc_loop_monitor_68 = new(upc_loop_intf_68,upc_loop_csv_dumper_68);
    upc_loop_csv_dumper_69 = new("./upc_loop_status69.csv");
    upc_loop_monitor_69 = new(upc_loop_intf_69,upc_loop_csv_dumper_69);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(module_monitor_53);
    sample_manager_inst.add_one_monitor(module_monitor_54);
    sample_manager_inst.add_one_monitor(module_monitor_55);
    sample_manager_inst.add_one_monitor(module_monitor_56);
    sample_manager_inst.add_one_monitor(module_monitor_57);
    sample_manager_inst.add_one_monitor(module_monitor_58);
    sample_manager_inst.add_one_monitor(module_monitor_59);
    sample_manager_inst.add_one_monitor(module_monitor_60);
    sample_manager_inst.add_one_monitor(module_monitor_61);
    sample_manager_inst.add_one_monitor(module_monitor_62);
    sample_manager_inst.add_one_monitor(module_monitor_63);
    sample_manager_inst.add_one_monitor(module_monitor_64);
    sample_manager_inst.add_one_monitor(module_monitor_65);
    sample_manager_inst.add_one_monitor(module_monitor_66);
    sample_manager_inst.add_one_monitor(module_monitor_67);
    sample_manager_inst.add_one_monitor(module_monitor_68);
    sample_manager_inst.add_one_monitor(module_monitor_69);
    sample_manager_inst.add_one_monitor(module_monitor_70);
    sample_manager_inst.add_one_monitor(module_monitor_71);
    sample_manager_inst.add_one_monitor(module_monitor_72);
    sample_manager_inst.add_one_monitor(module_monitor_73);
    sample_manager_inst.add_one_monitor(module_monitor_74);
    sample_manager_inst.add_one_monitor(module_monitor_75);
    sample_manager_inst.add_one_monitor(module_monitor_76);
    sample_manager_inst.add_one_monitor(module_monitor_77);
    sample_manager_inst.add_one_monitor(module_monitor_78);
    sample_manager_inst.add_one_monitor(module_monitor_79);
    sample_manager_inst.add_one_monitor(module_monitor_80);
    sample_manager_inst.add_one_monitor(module_monitor_81);
    sample_manager_inst.add_one_monitor(module_monitor_82);
    sample_manager_inst.add_one_monitor(module_monitor_83);
    sample_manager_inst.add_one_monitor(module_monitor_84);
    sample_manager_inst.add_one_monitor(module_monitor_85);
    sample_manager_inst.add_one_monitor(module_monitor_86);
    sample_manager_inst.add_one_monitor(module_monitor_87);
    sample_manager_inst.add_one_monitor(module_monitor_88);
    sample_manager_inst.add_one_monitor(module_monitor_89);
    sample_manager_inst.add_one_monitor(module_monitor_90);
    sample_manager_inst.add_one_monitor(module_monitor_91);
    sample_manager_inst.add_one_monitor(module_monitor_92);
    sample_manager_inst.add_one_monitor(module_monitor_93);
    sample_manager_inst.add_one_monitor(module_monitor_94);
    sample_manager_inst.add_one_monitor(module_monitor_95);
    sample_manager_inst.add_one_monitor(module_monitor_96);
    sample_manager_inst.add_one_monitor(module_monitor_97);
    sample_manager_inst.add_one_monitor(module_monitor_98);
    sample_manager_inst.add_one_monitor(module_monitor_99);
    sample_manager_inst.add_one_monitor(module_monitor_100);
    sample_manager_inst.add_one_monitor(module_monitor_101);
    sample_manager_inst.add_one_monitor(module_monitor_102);
    sample_manager_inst.add_one_monitor(module_monitor_103);
    sample_manager_inst.add_one_monitor(module_monitor_104);
    sample_manager_inst.add_one_monitor(module_monitor_105);
    sample_manager_inst.add_one_monitor(module_monitor_106);
    sample_manager_inst.add_one_monitor(module_monitor_107);
    sample_manager_inst.add_one_monitor(module_monitor_108);
    sample_manager_inst.add_one_monitor(module_monitor_109);
    sample_manager_inst.add_one_monitor(module_monitor_110);
    sample_manager_inst.add_one_monitor(module_monitor_111);
    sample_manager_inst.add_one_monitor(module_monitor_112);
    sample_manager_inst.add_one_monitor(module_monitor_113);
    sample_manager_inst.add_one_monitor(module_monitor_114);
    sample_manager_inst.add_one_monitor(module_monitor_115);
    sample_manager_inst.add_one_monitor(module_monitor_116);
    sample_manager_inst.add_one_monitor(module_monitor_117);
    sample_manager_inst.add_one_monitor(module_monitor_118);
    sample_manager_inst.add_one_monitor(module_monitor_119);
    sample_manager_inst.add_one_monitor(module_monitor_120);
    sample_manager_inst.add_one_monitor(module_monitor_121);
    sample_manager_inst.add_one_monitor(module_monitor_122);
    sample_manager_inst.add_one_monitor(module_monitor_123);
    sample_manager_inst.add_one_monitor(module_monitor_124);
    sample_manager_inst.add_one_monitor(module_monitor_125);
    sample_manager_inst.add_one_monitor(module_monitor_126);
    sample_manager_inst.add_one_monitor(module_monitor_127);
    sample_manager_inst.add_one_monitor(module_monitor_128);
    sample_manager_inst.add_one_monitor(module_monitor_129);
    sample_manager_inst.add_one_monitor(module_monitor_130);
    sample_manager_inst.add_one_monitor(module_monitor_131);
    sample_manager_inst.add_one_monitor(module_monitor_132);
    sample_manager_inst.add_one_monitor(module_monitor_133);
    sample_manager_inst.add_one_monitor(module_monitor_134);
    sample_manager_inst.add_one_monitor(module_monitor_135);
    sample_manager_inst.add_one_monitor(module_monitor_136);
    sample_manager_inst.add_one_monitor(module_monitor_137);
    sample_manager_inst.add_one_monitor(module_monitor_138);
    sample_manager_inst.add_one_monitor(module_monitor_139);
    sample_manager_inst.add_one_monitor(module_monitor_140);
    sample_manager_inst.add_one_monitor(module_monitor_141);
    sample_manager_inst.add_one_monitor(module_monitor_142);
    sample_manager_inst.add_one_monitor(module_monitor_143);
    sample_manager_inst.add_one_monitor(module_monitor_144);
    sample_manager_inst.add_one_monitor(module_monitor_145);
    sample_manager_inst.add_one_monitor(module_monitor_146);
    sample_manager_inst.add_one_monitor(module_monitor_147);
    sample_manager_inst.add_one_monitor(module_monitor_148);
    sample_manager_inst.add_one_monitor(module_monitor_149);
    sample_manager_inst.add_one_monitor(module_monitor_150);
    sample_manager_inst.add_one_monitor(module_monitor_151);
    sample_manager_inst.add_one_monitor(module_monitor_152);
    sample_manager_inst.add_one_monitor(module_monitor_153);
    sample_manager_inst.add_one_monitor(module_monitor_154);
    sample_manager_inst.add_one_monitor(module_monitor_155);
    sample_manager_inst.add_one_monitor(module_monitor_156);
    sample_manager_inst.add_one_monitor(module_monitor_157);
    sample_manager_inst.add_one_monitor(module_monitor_158);
    sample_manager_inst.add_one_monitor(module_monitor_159);
    sample_manager_inst.add_one_monitor(module_monitor_160);
    sample_manager_inst.add_one_monitor(module_monitor_161);
    sample_manager_inst.add_one_monitor(module_monitor_162);
    sample_manager_inst.add_one_monitor(module_monitor_163);
    sample_manager_inst.add_one_monitor(module_monitor_164);
    sample_manager_inst.add_one_monitor(module_monitor_165);
    sample_manager_inst.add_one_monitor(module_monitor_166);
    sample_manager_inst.add_one_monitor(module_monitor_167);
    sample_manager_inst.add_one_monitor(module_monitor_168);
    sample_manager_inst.add_one_monitor(module_monitor_169);
    sample_manager_inst.add_one_monitor(module_monitor_170);
    sample_manager_inst.add_one_monitor(module_monitor_171);
    sample_manager_inst.add_one_monitor(module_monitor_172);
    sample_manager_inst.add_one_monitor(module_monitor_173);
    sample_manager_inst.add_one_monitor(module_monitor_174);
    sample_manager_inst.add_one_monitor(module_monitor_175);
    sample_manager_inst.add_one_monitor(module_monitor_176);
    sample_manager_inst.add_one_monitor(module_monitor_177);
    sample_manager_inst.add_one_monitor(module_monitor_178);
    sample_manager_inst.add_one_monitor(module_monitor_179);
    sample_manager_inst.add_one_monitor(module_monitor_180);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_1);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_2);
    sample_manager_inst.add_one_monitor(pp_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_10);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_11);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_12);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_13);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_14);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_15);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_16);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_17);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_18);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_19);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_20);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_21);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_22);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_23);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_24);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_25);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_26);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_27);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_28);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_29);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_30);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_31);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_32);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_33);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_34);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_2);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_3);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_4);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_5);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_6);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_7);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_8);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_9);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_10);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_11);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_12);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_13);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_14);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_15);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_16);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_17);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_18);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_19);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_20);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_21);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_22);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_23);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_24);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_25);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_26);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_27);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_28);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_29);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_30);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_31);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_32);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_33);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_34);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_35);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_36);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_37);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_38);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_39);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_40);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_41);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_42);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_43);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_44);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_45);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_46);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_47);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_48);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_49);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_50);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_51);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_52);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_53);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_54);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_55);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_56);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_57);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_58);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_59);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_60);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_61);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_62);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_63);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_64);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_65);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_66);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_67);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_68);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_69);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
