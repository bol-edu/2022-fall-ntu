// initial a empty file
