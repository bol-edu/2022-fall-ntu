defparam AESL_inst_example.data_channel1_U.DEPTH = 'd11;
defparam AESL_inst_example.data_channel1_U.ADDR_WIDTH = 'd4;
defparam AESL_inst_example.data_channel2_U.DEPTH = 'd2;
defparam AESL_inst_example.data_channel2_U.ADDR_WIDTH = 'd1;
defparam AESL_inst_example.proc_1_U0.data_channel1_U.DEPTH = 'd11;
defparam AESL_inst_example.proc_1_U0.data_channel1_U.ADDR_WIDTH = 'd4;
defparam AESL_inst_example.proc_1_U0.data_channel2_U.DEPTH = 'd4;
defparam AESL_inst_example.proc_1_U0.data_channel2_U.ADDR_WIDTH = 'd2;
defparam AESL_inst_example.proc_2_U0.data_channel1_U.DEPTH = 'd11;
defparam AESL_inst_example.proc_2_U0.data_channel1_U.ADDR_WIDTH = 'd4;
defparam AESL_inst_example.proc_2_U0.data_channel2_U.DEPTH = 'd2;
defparam AESL_inst_example.proc_2_U0.data_channel2_U.ADDR_WIDTH = 'd1;
