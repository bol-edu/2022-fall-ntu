defparam AESL_inst_canny.upperThresh_c_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.upperThresh_c_U.ADDR_WIDTH = 32'd10;
defparam AESL_inst_canny.lowerThresh_c_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.lowerThresh_c_U.ADDR_WIDTH = 32'd10;
defparam AESL_inst_canny.x_sobel_V_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.x_sobel_V_U.ADDR_WIDTH = 32'd10;
defparam AESL_inst_canny.y_sobel_V_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.y_sobel_V_U.ADDR_WIDTH = 32'd10;
defparam AESL_inst_canny.y_sobel_7_V_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.y_sobel_7_V_U.ADDR_WIDTH = 32'd10;
defparam AESL_inst_canny.magnitude_V_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.magnitude_V_U.ADDR_WIDTH = 32'd10;
defparam AESL_inst_canny.tangent_y_V_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.tangent_y_V_U.ADDR_WIDTH = 32'd10;
defparam AESL_inst_canny.tangent_x_225_V_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.tangent_x_225_V_U.ADDR_WIDTH = 32'd10;
defparam AESL_inst_canny.tangent_x_675_V_U.DEPTH = 11'd1000;
defparam AESL_inst_canny.tangent_x_675_V_U.ADDR_WIDTH = 32'd10;
